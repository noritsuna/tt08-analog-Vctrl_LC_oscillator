VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_noritsuna_Vctrl_LC_oscillator
  CLASS BLOCK ;
  FOREIGN tt_um_noritsuna_Vctrl_LC_oscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN vout_p
    ANTENNAGATEAREA 2000.000000 ;
    ANTENNADIFFAREA 1094.500000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END vout_p
  PIN vout_n
    ANTENNAGATEAREA 2000.000000 ;
    ANTENNADIFFAREA 1094.500000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END vout_n
  PIN vctrl
    ANTENNADIFFAREA 35.171600 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END vctrl
  PIN ibias
    ANTENNAGATEAREA 50.000000 ;
    ANTENNADIFFAREA 12.500000 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ibias
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 47.455997 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    ANTENNAGATEAREA 2000.000000 ;
    ANTENNADIFFAREA 1094.500000 ;
    PORT
      LAYER met4 ;
        RECT 7.000 5.000 9.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER pwell ;
        RECT 118.850 172.350 142.570 172.840 ;
        RECT 118.850 119.610 119.340 172.350 ;
      LAYER nwell ;
        RECT 119.990 120.370 141.440 171.630 ;
      LAYER pwell ;
        RECT 142.080 119.610 142.570 172.350 ;
        RECT 118.850 119.120 142.570 119.610 ;
        RECT 11.700 108.870 117.880 114.900 ;
        RECT 11.700 107.700 12.260 108.870 ;
        RECT 117.320 107.700 117.880 108.870 ;
        RECT 11.700 95.520 117.880 107.700 ;
        RECT 11.700 94.350 12.260 95.520 ;
        RECT 117.320 94.350 117.880 95.520 ;
        RECT 11.700 82.170 117.880 94.350 ;
        RECT 11.700 81.000 12.260 82.170 ;
        RECT 117.320 81.000 117.880 82.170 ;
        RECT 11.700 68.820 117.880 81.000 ;
        RECT 11.700 67.650 12.260 68.820 ;
        RECT 117.320 67.650 117.880 68.820 ;
        RECT 11.700 61.620 117.880 67.650 ;
        RECT 52.000 4.870 75.750 12.010 ;
      LAYER li1 ;
        RECT 118.980 172.480 142.440 172.710 ;
        RECT 118.980 119.480 119.210 172.480 ;
        RECT 120.830 171.230 140.600 171.400 ;
        RECT 120.260 121.170 120.430 170.820 ;
        RECT 141.000 121.170 141.170 170.820 ;
        RECT 120.830 120.600 140.600 120.770 ;
        RECT 142.210 119.480 142.440 172.480 ;
        RECT 118.980 119.250 142.440 119.480 ;
        RECT 11.830 114.470 117.750 114.770 ;
        RECT 11.830 102.100 12.130 114.470 ;
        RECT 12.640 109.170 12.810 113.820 ;
        RECT 13.540 109.170 13.710 113.820 ;
        RECT 14.540 109.170 14.710 113.820 ;
        RECT 15.540 109.170 15.710 113.820 ;
        RECT 16.540 109.170 16.710 113.820 ;
        RECT 17.540 109.170 17.710 113.820 ;
        RECT 18.540 109.170 18.710 113.820 ;
        RECT 19.540 109.170 19.710 113.820 ;
        RECT 20.540 109.170 20.710 113.820 ;
        RECT 21.540 109.170 21.710 113.820 ;
        RECT 22.440 109.170 22.610 113.820 ;
        RECT 23.120 109.170 23.290 113.820 ;
        RECT 24.020 109.170 24.190 113.820 ;
        RECT 25.020 109.170 25.190 113.820 ;
        RECT 26.020 109.170 26.190 113.820 ;
        RECT 27.020 109.170 27.190 113.820 ;
        RECT 28.020 109.170 28.190 113.820 ;
        RECT 29.020 109.170 29.190 113.820 ;
        RECT 30.020 109.170 30.190 113.820 ;
        RECT 31.020 109.170 31.190 113.820 ;
        RECT 32.020 109.170 32.190 113.820 ;
        RECT 32.920 109.170 33.090 113.820 ;
        RECT 33.600 109.170 33.770 113.820 ;
        RECT 34.500 109.170 34.670 113.820 ;
        RECT 35.500 109.170 35.670 113.820 ;
        RECT 36.500 109.170 36.670 113.820 ;
        RECT 37.500 109.170 37.670 113.820 ;
        RECT 38.500 109.170 38.670 113.820 ;
        RECT 39.500 109.170 39.670 113.820 ;
        RECT 40.500 109.170 40.670 113.820 ;
        RECT 41.500 109.170 41.670 113.820 ;
        RECT 42.500 109.170 42.670 113.820 ;
        RECT 43.400 109.170 43.570 113.820 ;
        RECT 44.080 109.170 44.250 113.820 ;
        RECT 44.980 109.170 45.150 113.820 ;
        RECT 45.980 109.170 46.150 113.820 ;
        RECT 46.980 109.170 47.150 113.820 ;
        RECT 47.980 109.170 48.150 113.820 ;
        RECT 48.980 109.170 49.150 113.820 ;
        RECT 49.980 109.170 50.150 113.820 ;
        RECT 50.980 109.170 51.150 113.820 ;
        RECT 51.980 109.170 52.150 113.820 ;
        RECT 52.980 109.170 53.150 113.820 ;
        RECT 53.880 109.170 54.050 113.820 ;
        RECT 54.560 109.170 54.730 113.820 ;
        RECT 55.460 109.170 55.630 113.820 ;
        RECT 56.460 109.170 56.630 113.820 ;
        RECT 57.460 109.170 57.630 113.820 ;
        RECT 58.460 109.170 58.630 113.820 ;
        RECT 59.460 109.170 59.630 113.820 ;
        RECT 60.460 109.170 60.630 113.820 ;
        RECT 61.460 109.170 61.630 113.820 ;
        RECT 62.460 109.170 62.630 113.820 ;
        RECT 63.460 109.170 63.630 113.820 ;
        RECT 64.360 109.170 64.530 113.820 ;
        RECT 65.040 109.170 65.210 113.820 ;
        RECT 65.940 109.170 66.110 113.820 ;
        RECT 66.940 109.170 67.110 113.820 ;
        RECT 67.940 109.170 68.110 113.820 ;
        RECT 68.940 109.170 69.110 113.820 ;
        RECT 69.940 109.170 70.110 113.820 ;
        RECT 70.940 109.170 71.110 113.820 ;
        RECT 71.940 109.170 72.110 113.820 ;
        RECT 72.940 109.170 73.110 113.820 ;
        RECT 73.940 109.170 74.110 113.820 ;
        RECT 74.840 109.170 75.010 113.820 ;
        RECT 75.520 109.170 75.690 113.820 ;
        RECT 76.420 109.170 76.590 113.820 ;
        RECT 77.420 109.170 77.590 113.820 ;
        RECT 78.420 109.170 78.590 113.820 ;
        RECT 79.420 109.170 79.590 113.820 ;
        RECT 80.420 109.170 80.590 113.820 ;
        RECT 81.420 109.170 81.590 113.820 ;
        RECT 82.420 109.170 82.590 113.820 ;
        RECT 83.420 109.170 83.590 113.820 ;
        RECT 84.420 109.170 84.590 113.820 ;
        RECT 85.320 109.170 85.490 113.820 ;
        RECT 86.000 109.170 86.170 113.820 ;
        RECT 86.900 109.170 87.070 113.820 ;
        RECT 87.900 109.170 88.070 113.820 ;
        RECT 88.900 109.170 89.070 113.820 ;
        RECT 89.900 109.170 90.070 113.820 ;
        RECT 90.900 109.170 91.070 113.820 ;
        RECT 91.900 109.170 92.070 113.820 ;
        RECT 92.900 109.170 93.070 113.820 ;
        RECT 93.900 109.170 94.070 113.820 ;
        RECT 94.900 109.170 95.070 113.820 ;
        RECT 95.800 109.170 95.970 113.820 ;
        RECT 96.480 109.170 96.650 113.820 ;
        RECT 97.380 109.170 97.550 113.820 ;
        RECT 98.380 109.170 98.550 113.820 ;
        RECT 99.380 109.170 99.550 113.820 ;
        RECT 100.380 109.170 100.550 113.820 ;
        RECT 101.380 109.170 101.550 113.820 ;
        RECT 102.380 109.170 102.550 113.820 ;
        RECT 103.380 109.170 103.550 113.820 ;
        RECT 104.380 109.170 104.550 113.820 ;
        RECT 105.380 109.170 105.550 113.820 ;
        RECT 106.280 109.170 106.450 113.820 ;
        RECT 106.960 109.170 107.130 113.820 ;
        RECT 107.860 109.170 108.030 113.820 ;
        RECT 108.860 109.170 109.030 113.820 ;
        RECT 109.860 109.170 110.030 113.820 ;
        RECT 110.860 109.170 111.030 113.820 ;
        RECT 111.860 109.170 112.030 113.820 ;
        RECT 112.860 109.170 113.030 113.820 ;
        RECT 113.860 109.170 114.030 113.820 ;
        RECT 114.860 109.170 115.030 113.820 ;
        RECT 115.860 109.170 116.030 113.820 ;
        RECT 116.760 109.170 116.930 113.820 ;
        RECT 12.960 108.540 13.290 108.710 ;
        RECT 13.960 108.540 14.290 108.710 ;
        RECT 14.960 108.540 15.290 108.710 ;
        RECT 15.960 108.540 16.290 108.710 ;
        RECT 16.960 108.540 17.290 108.710 ;
        RECT 17.960 108.540 18.290 108.710 ;
        RECT 18.960 108.540 19.290 108.710 ;
        RECT 19.960 108.540 20.290 108.710 ;
        RECT 20.960 108.540 21.290 108.710 ;
        RECT 21.960 108.540 22.290 108.710 ;
        RECT 23.440 108.540 23.770 108.710 ;
        RECT 24.440 108.540 24.770 108.710 ;
        RECT 25.440 108.540 25.770 108.710 ;
        RECT 26.440 108.540 26.770 108.710 ;
        RECT 27.440 108.540 27.770 108.710 ;
        RECT 28.440 108.540 28.770 108.710 ;
        RECT 29.440 108.540 29.770 108.710 ;
        RECT 30.440 108.540 30.770 108.710 ;
        RECT 31.440 108.540 31.770 108.710 ;
        RECT 32.440 108.540 32.770 108.710 ;
        RECT 33.920 108.540 34.250 108.710 ;
        RECT 34.920 108.540 35.250 108.710 ;
        RECT 35.920 108.540 36.250 108.710 ;
        RECT 36.920 108.540 37.250 108.710 ;
        RECT 37.920 108.540 38.250 108.710 ;
        RECT 38.920 108.540 39.250 108.710 ;
        RECT 39.920 108.540 40.250 108.710 ;
        RECT 40.920 108.540 41.250 108.710 ;
        RECT 41.920 108.540 42.250 108.710 ;
        RECT 42.920 108.540 43.250 108.710 ;
        RECT 44.400 108.540 44.730 108.710 ;
        RECT 45.400 108.540 45.730 108.710 ;
        RECT 46.400 108.540 46.730 108.710 ;
        RECT 47.400 108.540 47.730 108.710 ;
        RECT 48.400 108.540 48.730 108.710 ;
        RECT 49.400 108.540 49.730 108.710 ;
        RECT 50.400 108.540 50.730 108.710 ;
        RECT 51.400 108.540 51.730 108.710 ;
        RECT 52.400 108.540 52.730 108.710 ;
        RECT 53.400 108.540 53.730 108.710 ;
        RECT 54.880 108.540 55.210 108.710 ;
        RECT 55.880 108.540 56.210 108.710 ;
        RECT 56.880 108.540 57.210 108.710 ;
        RECT 57.880 108.540 58.210 108.710 ;
        RECT 58.880 108.540 59.210 108.710 ;
        RECT 59.880 108.540 60.210 108.710 ;
        RECT 60.880 108.540 61.210 108.710 ;
        RECT 61.880 108.540 62.210 108.710 ;
        RECT 62.880 108.540 63.210 108.710 ;
        RECT 63.880 108.540 64.210 108.710 ;
        RECT 65.360 108.540 65.690 108.710 ;
        RECT 66.360 108.540 66.690 108.710 ;
        RECT 67.360 108.540 67.690 108.710 ;
        RECT 68.360 108.540 68.690 108.710 ;
        RECT 69.360 108.540 69.690 108.710 ;
        RECT 70.360 108.540 70.690 108.710 ;
        RECT 71.360 108.540 71.690 108.710 ;
        RECT 72.360 108.540 72.690 108.710 ;
        RECT 73.360 108.540 73.690 108.710 ;
        RECT 74.360 108.540 74.690 108.710 ;
        RECT 75.840 108.540 76.170 108.710 ;
        RECT 76.840 108.540 77.170 108.710 ;
        RECT 77.840 108.540 78.170 108.710 ;
        RECT 78.840 108.540 79.170 108.710 ;
        RECT 79.840 108.540 80.170 108.710 ;
        RECT 80.840 108.540 81.170 108.710 ;
        RECT 81.840 108.540 82.170 108.710 ;
        RECT 82.840 108.540 83.170 108.710 ;
        RECT 83.840 108.540 84.170 108.710 ;
        RECT 84.840 108.540 85.170 108.710 ;
        RECT 86.320 108.540 86.650 108.710 ;
        RECT 87.320 108.540 87.650 108.710 ;
        RECT 88.320 108.540 88.650 108.710 ;
        RECT 89.320 108.540 89.650 108.710 ;
        RECT 90.320 108.540 90.650 108.710 ;
        RECT 91.320 108.540 91.650 108.710 ;
        RECT 92.320 108.540 92.650 108.710 ;
        RECT 93.320 108.540 93.650 108.710 ;
        RECT 94.320 108.540 94.650 108.710 ;
        RECT 95.320 108.540 95.650 108.710 ;
        RECT 96.800 108.540 97.130 108.710 ;
        RECT 97.800 108.540 98.130 108.710 ;
        RECT 98.800 108.540 99.130 108.710 ;
        RECT 99.800 108.540 100.130 108.710 ;
        RECT 100.800 108.540 101.130 108.710 ;
        RECT 101.800 108.540 102.130 108.710 ;
        RECT 102.800 108.540 103.130 108.710 ;
        RECT 103.800 108.540 104.130 108.710 ;
        RECT 104.800 108.540 105.130 108.710 ;
        RECT 105.800 108.540 106.130 108.710 ;
        RECT 107.280 108.540 107.610 108.710 ;
        RECT 108.280 108.540 108.610 108.710 ;
        RECT 109.280 108.540 109.610 108.710 ;
        RECT 110.280 108.540 110.610 108.710 ;
        RECT 111.280 108.540 111.610 108.710 ;
        RECT 112.280 108.540 112.610 108.710 ;
        RECT 113.280 108.540 113.610 108.710 ;
        RECT 114.280 108.540 114.610 108.710 ;
        RECT 115.280 108.540 115.610 108.710 ;
        RECT 116.280 108.540 116.610 108.710 ;
        RECT 12.970 107.860 13.300 108.030 ;
        RECT 13.970 107.860 14.300 108.030 ;
        RECT 14.970 107.860 15.300 108.030 ;
        RECT 15.970 107.860 16.300 108.030 ;
        RECT 16.970 107.860 17.300 108.030 ;
        RECT 17.970 107.860 18.300 108.030 ;
        RECT 18.970 107.860 19.300 108.030 ;
        RECT 19.970 107.860 20.300 108.030 ;
        RECT 20.970 107.860 21.300 108.030 ;
        RECT 21.970 107.860 22.300 108.030 ;
        RECT 23.450 107.860 23.780 108.030 ;
        RECT 24.450 107.860 24.780 108.030 ;
        RECT 25.450 107.860 25.780 108.030 ;
        RECT 26.450 107.860 26.780 108.030 ;
        RECT 27.450 107.860 27.780 108.030 ;
        RECT 28.450 107.860 28.780 108.030 ;
        RECT 29.450 107.860 29.780 108.030 ;
        RECT 30.450 107.860 30.780 108.030 ;
        RECT 31.450 107.860 31.780 108.030 ;
        RECT 32.450 107.860 32.780 108.030 ;
        RECT 33.930 107.860 34.260 108.030 ;
        RECT 34.930 107.860 35.260 108.030 ;
        RECT 35.930 107.860 36.260 108.030 ;
        RECT 36.930 107.860 37.260 108.030 ;
        RECT 37.930 107.860 38.260 108.030 ;
        RECT 38.930 107.860 39.260 108.030 ;
        RECT 39.930 107.860 40.260 108.030 ;
        RECT 40.930 107.860 41.260 108.030 ;
        RECT 41.930 107.860 42.260 108.030 ;
        RECT 42.930 107.860 43.260 108.030 ;
        RECT 44.410 107.860 44.740 108.030 ;
        RECT 45.410 107.860 45.740 108.030 ;
        RECT 46.410 107.860 46.740 108.030 ;
        RECT 47.410 107.860 47.740 108.030 ;
        RECT 48.410 107.860 48.740 108.030 ;
        RECT 49.410 107.860 49.740 108.030 ;
        RECT 50.410 107.860 50.740 108.030 ;
        RECT 51.410 107.860 51.740 108.030 ;
        RECT 52.410 107.860 52.740 108.030 ;
        RECT 53.410 107.860 53.740 108.030 ;
        RECT 54.890 107.860 55.220 108.030 ;
        RECT 55.890 107.860 56.220 108.030 ;
        RECT 56.890 107.860 57.220 108.030 ;
        RECT 57.890 107.860 58.220 108.030 ;
        RECT 58.890 107.860 59.220 108.030 ;
        RECT 59.890 107.860 60.220 108.030 ;
        RECT 60.890 107.860 61.220 108.030 ;
        RECT 61.890 107.860 62.220 108.030 ;
        RECT 62.890 107.860 63.220 108.030 ;
        RECT 63.890 107.860 64.220 108.030 ;
        RECT 65.370 107.860 65.700 108.030 ;
        RECT 66.370 107.860 66.700 108.030 ;
        RECT 67.370 107.860 67.700 108.030 ;
        RECT 68.370 107.860 68.700 108.030 ;
        RECT 69.370 107.860 69.700 108.030 ;
        RECT 70.370 107.860 70.700 108.030 ;
        RECT 71.370 107.860 71.700 108.030 ;
        RECT 72.370 107.860 72.700 108.030 ;
        RECT 73.370 107.860 73.700 108.030 ;
        RECT 74.370 107.860 74.700 108.030 ;
        RECT 75.850 107.860 76.180 108.030 ;
        RECT 76.850 107.860 77.180 108.030 ;
        RECT 77.850 107.860 78.180 108.030 ;
        RECT 78.850 107.860 79.180 108.030 ;
        RECT 79.850 107.860 80.180 108.030 ;
        RECT 80.850 107.860 81.180 108.030 ;
        RECT 81.850 107.860 82.180 108.030 ;
        RECT 82.850 107.860 83.180 108.030 ;
        RECT 83.850 107.860 84.180 108.030 ;
        RECT 84.850 107.860 85.180 108.030 ;
        RECT 86.330 107.860 86.660 108.030 ;
        RECT 87.330 107.860 87.660 108.030 ;
        RECT 88.330 107.860 88.660 108.030 ;
        RECT 89.330 107.860 89.660 108.030 ;
        RECT 90.330 107.860 90.660 108.030 ;
        RECT 91.330 107.860 91.660 108.030 ;
        RECT 92.330 107.860 92.660 108.030 ;
        RECT 93.330 107.860 93.660 108.030 ;
        RECT 94.330 107.860 94.660 108.030 ;
        RECT 95.330 107.860 95.660 108.030 ;
        RECT 96.810 107.860 97.140 108.030 ;
        RECT 97.810 107.860 98.140 108.030 ;
        RECT 98.810 107.860 99.140 108.030 ;
        RECT 99.810 107.860 100.140 108.030 ;
        RECT 100.810 107.860 101.140 108.030 ;
        RECT 101.810 107.860 102.140 108.030 ;
        RECT 102.810 107.860 103.140 108.030 ;
        RECT 103.810 107.860 104.140 108.030 ;
        RECT 104.810 107.860 105.140 108.030 ;
        RECT 105.810 107.860 106.140 108.030 ;
        RECT 107.290 107.860 107.620 108.030 ;
        RECT 108.290 107.860 108.620 108.030 ;
        RECT 109.290 107.860 109.620 108.030 ;
        RECT 110.290 107.860 110.620 108.030 ;
        RECT 111.290 107.860 111.620 108.030 ;
        RECT 112.290 107.860 112.620 108.030 ;
        RECT 113.290 107.860 113.620 108.030 ;
        RECT 114.290 107.860 114.620 108.030 ;
        RECT 115.290 107.860 115.620 108.030 ;
        RECT 116.290 107.860 116.620 108.030 ;
        RECT 12.650 102.750 12.820 107.400 ;
        RECT 13.550 102.750 13.720 107.400 ;
        RECT 14.550 102.750 14.720 107.400 ;
        RECT 15.550 102.750 15.720 107.400 ;
        RECT 16.550 102.750 16.720 107.400 ;
        RECT 17.550 102.750 17.720 107.400 ;
        RECT 18.550 102.750 18.720 107.400 ;
        RECT 19.550 102.750 19.720 107.400 ;
        RECT 20.550 102.750 20.720 107.400 ;
        RECT 21.550 102.750 21.720 107.400 ;
        RECT 22.450 102.750 22.620 107.400 ;
        RECT 23.130 102.750 23.300 107.400 ;
        RECT 24.030 102.750 24.200 107.400 ;
        RECT 25.030 102.750 25.200 107.400 ;
        RECT 26.030 102.750 26.200 107.400 ;
        RECT 27.030 102.750 27.200 107.400 ;
        RECT 28.030 102.750 28.200 107.400 ;
        RECT 29.030 102.750 29.200 107.400 ;
        RECT 30.030 102.750 30.200 107.400 ;
        RECT 31.030 102.750 31.200 107.400 ;
        RECT 32.030 102.750 32.200 107.400 ;
        RECT 32.930 102.750 33.100 107.400 ;
        RECT 33.610 102.750 33.780 107.400 ;
        RECT 34.510 102.750 34.680 107.400 ;
        RECT 35.510 102.750 35.680 107.400 ;
        RECT 36.510 102.750 36.680 107.400 ;
        RECT 37.510 102.750 37.680 107.400 ;
        RECT 38.510 102.750 38.680 107.400 ;
        RECT 39.510 102.750 39.680 107.400 ;
        RECT 40.510 102.750 40.680 107.400 ;
        RECT 41.510 102.750 41.680 107.400 ;
        RECT 42.510 102.750 42.680 107.400 ;
        RECT 43.410 102.750 43.580 107.400 ;
        RECT 44.090 102.750 44.260 107.400 ;
        RECT 44.990 102.750 45.160 107.400 ;
        RECT 45.990 102.750 46.160 107.400 ;
        RECT 46.990 102.750 47.160 107.400 ;
        RECT 47.990 102.750 48.160 107.400 ;
        RECT 48.990 102.750 49.160 107.400 ;
        RECT 49.990 102.750 50.160 107.400 ;
        RECT 50.990 102.750 51.160 107.400 ;
        RECT 51.990 102.750 52.160 107.400 ;
        RECT 52.990 102.750 53.160 107.400 ;
        RECT 53.890 102.750 54.060 107.400 ;
        RECT 54.570 102.750 54.740 107.400 ;
        RECT 55.470 102.750 55.640 107.400 ;
        RECT 56.470 102.750 56.640 107.400 ;
        RECT 57.470 102.750 57.640 107.400 ;
        RECT 58.470 102.750 58.640 107.400 ;
        RECT 59.470 102.750 59.640 107.400 ;
        RECT 60.470 102.750 60.640 107.400 ;
        RECT 61.470 102.750 61.640 107.400 ;
        RECT 62.470 102.750 62.640 107.400 ;
        RECT 63.470 102.750 63.640 107.400 ;
        RECT 64.370 102.750 64.540 107.400 ;
        RECT 65.050 102.750 65.220 107.400 ;
        RECT 65.950 102.750 66.120 107.400 ;
        RECT 66.950 102.750 67.120 107.400 ;
        RECT 67.950 102.750 68.120 107.400 ;
        RECT 68.950 102.750 69.120 107.400 ;
        RECT 69.950 102.750 70.120 107.400 ;
        RECT 70.950 102.750 71.120 107.400 ;
        RECT 71.950 102.750 72.120 107.400 ;
        RECT 72.950 102.750 73.120 107.400 ;
        RECT 73.950 102.750 74.120 107.400 ;
        RECT 74.850 102.750 75.020 107.400 ;
        RECT 75.530 102.750 75.700 107.400 ;
        RECT 76.430 102.750 76.600 107.400 ;
        RECT 77.430 102.750 77.600 107.400 ;
        RECT 78.430 102.750 78.600 107.400 ;
        RECT 79.430 102.750 79.600 107.400 ;
        RECT 80.430 102.750 80.600 107.400 ;
        RECT 81.430 102.750 81.600 107.400 ;
        RECT 82.430 102.750 82.600 107.400 ;
        RECT 83.430 102.750 83.600 107.400 ;
        RECT 84.430 102.750 84.600 107.400 ;
        RECT 85.330 102.750 85.500 107.400 ;
        RECT 86.010 102.750 86.180 107.400 ;
        RECT 86.910 102.750 87.080 107.400 ;
        RECT 87.910 102.750 88.080 107.400 ;
        RECT 88.910 102.750 89.080 107.400 ;
        RECT 89.910 102.750 90.080 107.400 ;
        RECT 90.910 102.750 91.080 107.400 ;
        RECT 91.910 102.750 92.080 107.400 ;
        RECT 92.910 102.750 93.080 107.400 ;
        RECT 93.910 102.750 94.080 107.400 ;
        RECT 94.910 102.750 95.080 107.400 ;
        RECT 95.810 102.750 95.980 107.400 ;
        RECT 96.490 102.750 96.660 107.400 ;
        RECT 97.390 102.750 97.560 107.400 ;
        RECT 98.390 102.750 98.560 107.400 ;
        RECT 99.390 102.750 99.560 107.400 ;
        RECT 100.390 102.750 100.560 107.400 ;
        RECT 101.390 102.750 101.560 107.400 ;
        RECT 102.390 102.750 102.560 107.400 ;
        RECT 103.390 102.750 103.560 107.400 ;
        RECT 104.390 102.750 104.560 107.400 ;
        RECT 105.390 102.750 105.560 107.400 ;
        RECT 106.290 102.750 106.460 107.400 ;
        RECT 106.970 102.750 107.140 107.400 ;
        RECT 107.870 102.750 108.040 107.400 ;
        RECT 108.870 102.750 109.040 107.400 ;
        RECT 109.870 102.750 110.040 107.400 ;
        RECT 110.870 102.750 111.040 107.400 ;
        RECT 111.870 102.750 112.040 107.400 ;
        RECT 112.870 102.750 113.040 107.400 ;
        RECT 113.870 102.750 114.040 107.400 ;
        RECT 114.870 102.750 115.040 107.400 ;
        RECT 115.870 102.750 116.040 107.400 ;
        RECT 116.770 102.750 116.940 107.400 ;
        RECT 117.450 102.100 117.750 114.470 ;
        RECT 11.830 101.800 117.750 102.100 ;
        RECT 11.830 101.120 117.750 101.420 ;
        RECT 11.830 88.750 12.130 101.120 ;
        RECT 12.640 95.820 12.810 100.470 ;
        RECT 13.540 95.820 13.710 100.470 ;
        RECT 14.540 95.820 14.710 100.470 ;
        RECT 15.540 95.820 15.710 100.470 ;
        RECT 16.540 95.820 16.710 100.470 ;
        RECT 17.540 95.820 17.710 100.470 ;
        RECT 18.540 95.820 18.710 100.470 ;
        RECT 19.540 95.820 19.710 100.470 ;
        RECT 20.540 95.820 20.710 100.470 ;
        RECT 21.540 95.820 21.710 100.470 ;
        RECT 22.440 95.820 22.610 100.470 ;
        RECT 23.120 95.820 23.290 100.470 ;
        RECT 24.020 95.820 24.190 100.470 ;
        RECT 25.020 95.820 25.190 100.470 ;
        RECT 26.020 95.820 26.190 100.470 ;
        RECT 27.020 95.820 27.190 100.470 ;
        RECT 28.020 95.820 28.190 100.470 ;
        RECT 29.020 95.820 29.190 100.470 ;
        RECT 30.020 95.820 30.190 100.470 ;
        RECT 31.020 95.820 31.190 100.470 ;
        RECT 32.020 95.820 32.190 100.470 ;
        RECT 32.920 95.820 33.090 100.470 ;
        RECT 33.600 95.820 33.770 100.470 ;
        RECT 34.500 95.820 34.670 100.470 ;
        RECT 35.500 95.820 35.670 100.470 ;
        RECT 36.500 95.820 36.670 100.470 ;
        RECT 37.500 95.820 37.670 100.470 ;
        RECT 38.500 95.820 38.670 100.470 ;
        RECT 39.500 95.820 39.670 100.470 ;
        RECT 40.500 95.820 40.670 100.470 ;
        RECT 41.500 95.820 41.670 100.470 ;
        RECT 42.500 95.820 42.670 100.470 ;
        RECT 43.400 95.820 43.570 100.470 ;
        RECT 44.080 95.820 44.250 100.470 ;
        RECT 44.980 95.820 45.150 100.470 ;
        RECT 45.980 95.820 46.150 100.470 ;
        RECT 46.980 95.820 47.150 100.470 ;
        RECT 47.980 95.820 48.150 100.470 ;
        RECT 48.980 95.820 49.150 100.470 ;
        RECT 49.980 95.820 50.150 100.470 ;
        RECT 50.980 95.820 51.150 100.470 ;
        RECT 51.980 95.820 52.150 100.470 ;
        RECT 52.980 95.820 53.150 100.470 ;
        RECT 53.880 95.820 54.050 100.470 ;
        RECT 54.560 95.820 54.730 100.470 ;
        RECT 55.460 95.820 55.630 100.470 ;
        RECT 56.460 95.820 56.630 100.470 ;
        RECT 57.460 95.820 57.630 100.470 ;
        RECT 58.460 95.820 58.630 100.470 ;
        RECT 59.460 95.820 59.630 100.470 ;
        RECT 60.460 95.820 60.630 100.470 ;
        RECT 61.460 95.820 61.630 100.470 ;
        RECT 62.460 95.820 62.630 100.470 ;
        RECT 63.460 95.820 63.630 100.470 ;
        RECT 64.360 95.820 64.530 100.470 ;
        RECT 65.040 95.820 65.210 100.470 ;
        RECT 65.940 95.820 66.110 100.470 ;
        RECT 66.940 95.820 67.110 100.470 ;
        RECT 67.940 95.820 68.110 100.470 ;
        RECT 68.940 95.820 69.110 100.470 ;
        RECT 69.940 95.820 70.110 100.470 ;
        RECT 70.940 95.820 71.110 100.470 ;
        RECT 71.940 95.820 72.110 100.470 ;
        RECT 72.940 95.820 73.110 100.470 ;
        RECT 73.940 95.820 74.110 100.470 ;
        RECT 74.840 95.820 75.010 100.470 ;
        RECT 75.520 95.820 75.690 100.470 ;
        RECT 76.420 95.820 76.590 100.470 ;
        RECT 77.420 95.820 77.590 100.470 ;
        RECT 78.420 95.820 78.590 100.470 ;
        RECT 79.420 95.820 79.590 100.470 ;
        RECT 80.420 95.820 80.590 100.470 ;
        RECT 81.420 95.820 81.590 100.470 ;
        RECT 82.420 95.820 82.590 100.470 ;
        RECT 83.420 95.820 83.590 100.470 ;
        RECT 84.420 95.820 84.590 100.470 ;
        RECT 85.320 95.820 85.490 100.470 ;
        RECT 86.000 95.820 86.170 100.470 ;
        RECT 86.900 95.820 87.070 100.470 ;
        RECT 87.900 95.820 88.070 100.470 ;
        RECT 88.900 95.820 89.070 100.470 ;
        RECT 89.900 95.820 90.070 100.470 ;
        RECT 90.900 95.820 91.070 100.470 ;
        RECT 91.900 95.820 92.070 100.470 ;
        RECT 92.900 95.820 93.070 100.470 ;
        RECT 93.900 95.820 94.070 100.470 ;
        RECT 94.900 95.820 95.070 100.470 ;
        RECT 95.800 95.820 95.970 100.470 ;
        RECT 96.480 95.820 96.650 100.470 ;
        RECT 97.380 95.820 97.550 100.470 ;
        RECT 98.380 95.820 98.550 100.470 ;
        RECT 99.380 95.820 99.550 100.470 ;
        RECT 100.380 95.820 100.550 100.470 ;
        RECT 101.380 95.820 101.550 100.470 ;
        RECT 102.380 95.820 102.550 100.470 ;
        RECT 103.380 95.820 103.550 100.470 ;
        RECT 104.380 95.820 104.550 100.470 ;
        RECT 105.380 95.820 105.550 100.470 ;
        RECT 106.280 95.820 106.450 100.470 ;
        RECT 106.960 95.820 107.130 100.470 ;
        RECT 107.860 95.820 108.030 100.470 ;
        RECT 108.860 95.820 109.030 100.470 ;
        RECT 109.860 95.820 110.030 100.470 ;
        RECT 110.860 95.820 111.030 100.470 ;
        RECT 111.860 95.820 112.030 100.470 ;
        RECT 112.860 95.820 113.030 100.470 ;
        RECT 113.860 95.820 114.030 100.470 ;
        RECT 114.860 95.820 115.030 100.470 ;
        RECT 115.860 95.820 116.030 100.470 ;
        RECT 116.760 95.820 116.930 100.470 ;
        RECT 12.960 95.190 13.290 95.360 ;
        RECT 13.960 95.190 14.290 95.360 ;
        RECT 14.960 95.190 15.290 95.360 ;
        RECT 15.960 95.190 16.290 95.360 ;
        RECT 16.960 95.190 17.290 95.360 ;
        RECT 17.960 95.190 18.290 95.360 ;
        RECT 18.960 95.190 19.290 95.360 ;
        RECT 19.960 95.190 20.290 95.360 ;
        RECT 20.960 95.190 21.290 95.360 ;
        RECT 21.960 95.190 22.290 95.360 ;
        RECT 23.440 95.190 23.770 95.360 ;
        RECT 24.440 95.190 24.770 95.360 ;
        RECT 25.440 95.190 25.770 95.360 ;
        RECT 26.440 95.190 26.770 95.360 ;
        RECT 27.440 95.190 27.770 95.360 ;
        RECT 28.440 95.190 28.770 95.360 ;
        RECT 29.440 95.190 29.770 95.360 ;
        RECT 30.440 95.190 30.770 95.360 ;
        RECT 31.440 95.190 31.770 95.360 ;
        RECT 32.440 95.190 32.770 95.360 ;
        RECT 33.920 95.190 34.250 95.360 ;
        RECT 34.920 95.190 35.250 95.360 ;
        RECT 35.920 95.190 36.250 95.360 ;
        RECT 36.920 95.190 37.250 95.360 ;
        RECT 37.920 95.190 38.250 95.360 ;
        RECT 38.920 95.190 39.250 95.360 ;
        RECT 39.920 95.190 40.250 95.360 ;
        RECT 40.920 95.190 41.250 95.360 ;
        RECT 41.920 95.190 42.250 95.360 ;
        RECT 42.920 95.190 43.250 95.360 ;
        RECT 44.400 95.190 44.730 95.360 ;
        RECT 45.400 95.190 45.730 95.360 ;
        RECT 46.400 95.190 46.730 95.360 ;
        RECT 47.400 95.190 47.730 95.360 ;
        RECT 48.400 95.190 48.730 95.360 ;
        RECT 49.400 95.190 49.730 95.360 ;
        RECT 50.400 95.190 50.730 95.360 ;
        RECT 51.400 95.190 51.730 95.360 ;
        RECT 52.400 95.190 52.730 95.360 ;
        RECT 53.400 95.190 53.730 95.360 ;
        RECT 54.880 95.190 55.210 95.360 ;
        RECT 55.880 95.190 56.210 95.360 ;
        RECT 56.880 95.190 57.210 95.360 ;
        RECT 57.880 95.190 58.210 95.360 ;
        RECT 58.880 95.190 59.210 95.360 ;
        RECT 59.880 95.190 60.210 95.360 ;
        RECT 60.880 95.190 61.210 95.360 ;
        RECT 61.880 95.190 62.210 95.360 ;
        RECT 62.880 95.190 63.210 95.360 ;
        RECT 63.880 95.190 64.210 95.360 ;
        RECT 65.360 95.190 65.690 95.360 ;
        RECT 66.360 95.190 66.690 95.360 ;
        RECT 67.360 95.190 67.690 95.360 ;
        RECT 68.360 95.190 68.690 95.360 ;
        RECT 69.360 95.190 69.690 95.360 ;
        RECT 70.360 95.190 70.690 95.360 ;
        RECT 71.360 95.190 71.690 95.360 ;
        RECT 72.360 95.190 72.690 95.360 ;
        RECT 73.360 95.190 73.690 95.360 ;
        RECT 74.360 95.190 74.690 95.360 ;
        RECT 75.840 95.190 76.170 95.360 ;
        RECT 76.840 95.190 77.170 95.360 ;
        RECT 77.840 95.190 78.170 95.360 ;
        RECT 78.840 95.190 79.170 95.360 ;
        RECT 79.840 95.190 80.170 95.360 ;
        RECT 80.840 95.190 81.170 95.360 ;
        RECT 81.840 95.190 82.170 95.360 ;
        RECT 82.840 95.190 83.170 95.360 ;
        RECT 83.840 95.190 84.170 95.360 ;
        RECT 84.840 95.190 85.170 95.360 ;
        RECT 86.320 95.190 86.650 95.360 ;
        RECT 87.320 95.190 87.650 95.360 ;
        RECT 88.320 95.190 88.650 95.360 ;
        RECT 89.320 95.190 89.650 95.360 ;
        RECT 90.320 95.190 90.650 95.360 ;
        RECT 91.320 95.190 91.650 95.360 ;
        RECT 92.320 95.190 92.650 95.360 ;
        RECT 93.320 95.190 93.650 95.360 ;
        RECT 94.320 95.190 94.650 95.360 ;
        RECT 95.320 95.190 95.650 95.360 ;
        RECT 96.800 95.190 97.130 95.360 ;
        RECT 97.800 95.190 98.130 95.360 ;
        RECT 98.800 95.190 99.130 95.360 ;
        RECT 99.800 95.190 100.130 95.360 ;
        RECT 100.800 95.190 101.130 95.360 ;
        RECT 101.800 95.190 102.130 95.360 ;
        RECT 102.800 95.190 103.130 95.360 ;
        RECT 103.800 95.190 104.130 95.360 ;
        RECT 104.800 95.190 105.130 95.360 ;
        RECT 105.800 95.190 106.130 95.360 ;
        RECT 107.280 95.190 107.610 95.360 ;
        RECT 108.280 95.190 108.610 95.360 ;
        RECT 109.280 95.190 109.610 95.360 ;
        RECT 110.280 95.190 110.610 95.360 ;
        RECT 111.280 95.190 111.610 95.360 ;
        RECT 112.280 95.190 112.610 95.360 ;
        RECT 113.280 95.190 113.610 95.360 ;
        RECT 114.280 95.190 114.610 95.360 ;
        RECT 115.280 95.190 115.610 95.360 ;
        RECT 116.280 95.190 116.610 95.360 ;
        RECT 12.970 94.510 13.300 94.680 ;
        RECT 13.970 94.510 14.300 94.680 ;
        RECT 14.970 94.510 15.300 94.680 ;
        RECT 15.970 94.510 16.300 94.680 ;
        RECT 16.970 94.510 17.300 94.680 ;
        RECT 17.970 94.510 18.300 94.680 ;
        RECT 18.970 94.510 19.300 94.680 ;
        RECT 19.970 94.510 20.300 94.680 ;
        RECT 20.970 94.510 21.300 94.680 ;
        RECT 21.970 94.510 22.300 94.680 ;
        RECT 23.450 94.510 23.780 94.680 ;
        RECT 24.450 94.510 24.780 94.680 ;
        RECT 25.450 94.510 25.780 94.680 ;
        RECT 26.450 94.510 26.780 94.680 ;
        RECT 27.450 94.510 27.780 94.680 ;
        RECT 28.450 94.510 28.780 94.680 ;
        RECT 29.450 94.510 29.780 94.680 ;
        RECT 30.450 94.510 30.780 94.680 ;
        RECT 31.450 94.510 31.780 94.680 ;
        RECT 32.450 94.510 32.780 94.680 ;
        RECT 33.930 94.510 34.260 94.680 ;
        RECT 34.930 94.510 35.260 94.680 ;
        RECT 35.930 94.510 36.260 94.680 ;
        RECT 36.930 94.510 37.260 94.680 ;
        RECT 37.930 94.510 38.260 94.680 ;
        RECT 38.930 94.510 39.260 94.680 ;
        RECT 39.930 94.510 40.260 94.680 ;
        RECT 40.930 94.510 41.260 94.680 ;
        RECT 41.930 94.510 42.260 94.680 ;
        RECT 42.930 94.510 43.260 94.680 ;
        RECT 44.410 94.510 44.740 94.680 ;
        RECT 45.410 94.510 45.740 94.680 ;
        RECT 46.410 94.510 46.740 94.680 ;
        RECT 47.410 94.510 47.740 94.680 ;
        RECT 48.410 94.510 48.740 94.680 ;
        RECT 49.410 94.510 49.740 94.680 ;
        RECT 50.410 94.510 50.740 94.680 ;
        RECT 51.410 94.510 51.740 94.680 ;
        RECT 52.410 94.510 52.740 94.680 ;
        RECT 53.410 94.510 53.740 94.680 ;
        RECT 54.890 94.510 55.220 94.680 ;
        RECT 55.890 94.510 56.220 94.680 ;
        RECT 56.890 94.510 57.220 94.680 ;
        RECT 57.890 94.510 58.220 94.680 ;
        RECT 58.890 94.510 59.220 94.680 ;
        RECT 59.890 94.510 60.220 94.680 ;
        RECT 60.890 94.510 61.220 94.680 ;
        RECT 61.890 94.510 62.220 94.680 ;
        RECT 62.890 94.510 63.220 94.680 ;
        RECT 63.890 94.510 64.220 94.680 ;
        RECT 65.370 94.510 65.700 94.680 ;
        RECT 66.370 94.510 66.700 94.680 ;
        RECT 67.370 94.510 67.700 94.680 ;
        RECT 68.370 94.510 68.700 94.680 ;
        RECT 69.370 94.510 69.700 94.680 ;
        RECT 70.370 94.510 70.700 94.680 ;
        RECT 71.370 94.510 71.700 94.680 ;
        RECT 72.370 94.510 72.700 94.680 ;
        RECT 73.370 94.510 73.700 94.680 ;
        RECT 74.370 94.510 74.700 94.680 ;
        RECT 75.850 94.510 76.180 94.680 ;
        RECT 76.850 94.510 77.180 94.680 ;
        RECT 77.850 94.510 78.180 94.680 ;
        RECT 78.850 94.510 79.180 94.680 ;
        RECT 79.850 94.510 80.180 94.680 ;
        RECT 80.850 94.510 81.180 94.680 ;
        RECT 81.850 94.510 82.180 94.680 ;
        RECT 82.850 94.510 83.180 94.680 ;
        RECT 83.850 94.510 84.180 94.680 ;
        RECT 84.850 94.510 85.180 94.680 ;
        RECT 86.330 94.510 86.660 94.680 ;
        RECT 87.330 94.510 87.660 94.680 ;
        RECT 88.330 94.510 88.660 94.680 ;
        RECT 89.330 94.510 89.660 94.680 ;
        RECT 90.330 94.510 90.660 94.680 ;
        RECT 91.330 94.510 91.660 94.680 ;
        RECT 92.330 94.510 92.660 94.680 ;
        RECT 93.330 94.510 93.660 94.680 ;
        RECT 94.330 94.510 94.660 94.680 ;
        RECT 95.330 94.510 95.660 94.680 ;
        RECT 96.810 94.510 97.140 94.680 ;
        RECT 97.810 94.510 98.140 94.680 ;
        RECT 98.810 94.510 99.140 94.680 ;
        RECT 99.810 94.510 100.140 94.680 ;
        RECT 100.810 94.510 101.140 94.680 ;
        RECT 101.810 94.510 102.140 94.680 ;
        RECT 102.810 94.510 103.140 94.680 ;
        RECT 103.810 94.510 104.140 94.680 ;
        RECT 104.810 94.510 105.140 94.680 ;
        RECT 105.810 94.510 106.140 94.680 ;
        RECT 107.290 94.510 107.620 94.680 ;
        RECT 108.290 94.510 108.620 94.680 ;
        RECT 109.290 94.510 109.620 94.680 ;
        RECT 110.290 94.510 110.620 94.680 ;
        RECT 111.290 94.510 111.620 94.680 ;
        RECT 112.290 94.510 112.620 94.680 ;
        RECT 113.290 94.510 113.620 94.680 ;
        RECT 114.290 94.510 114.620 94.680 ;
        RECT 115.290 94.510 115.620 94.680 ;
        RECT 116.290 94.510 116.620 94.680 ;
        RECT 12.650 89.400 12.820 94.050 ;
        RECT 13.550 89.400 13.720 94.050 ;
        RECT 14.550 89.400 14.720 94.050 ;
        RECT 15.550 89.400 15.720 94.050 ;
        RECT 16.550 89.400 16.720 94.050 ;
        RECT 17.550 89.400 17.720 94.050 ;
        RECT 18.550 89.400 18.720 94.050 ;
        RECT 19.550 89.400 19.720 94.050 ;
        RECT 20.550 89.400 20.720 94.050 ;
        RECT 21.550 89.400 21.720 94.050 ;
        RECT 22.450 89.400 22.620 94.050 ;
        RECT 23.130 89.400 23.300 94.050 ;
        RECT 24.030 89.400 24.200 94.050 ;
        RECT 25.030 89.400 25.200 94.050 ;
        RECT 26.030 89.400 26.200 94.050 ;
        RECT 27.030 89.400 27.200 94.050 ;
        RECT 28.030 89.400 28.200 94.050 ;
        RECT 29.030 89.400 29.200 94.050 ;
        RECT 30.030 89.400 30.200 94.050 ;
        RECT 31.030 89.400 31.200 94.050 ;
        RECT 32.030 89.400 32.200 94.050 ;
        RECT 32.930 89.400 33.100 94.050 ;
        RECT 33.610 89.400 33.780 94.050 ;
        RECT 34.510 89.400 34.680 94.050 ;
        RECT 35.510 89.400 35.680 94.050 ;
        RECT 36.510 89.400 36.680 94.050 ;
        RECT 37.510 89.400 37.680 94.050 ;
        RECT 38.510 89.400 38.680 94.050 ;
        RECT 39.510 89.400 39.680 94.050 ;
        RECT 40.510 89.400 40.680 94.050 ;
        RECT 41.510 89.400 41.680 94.050 ;
        RECT 42.510 89.400 42.680 94.050 ;
        RECT 43.410 89.400 43.580 94.050 ;
        RECT 44.090 89.400 44.260 94.050 ;
        RECT 44.990 89.400 45.160 94.050 ;
        RECT 45.990 89.400 46.160 94.050 ;
        RECT 46.990 89.400 47.160 94.050 ;
        RECT 47.990 89.400 48.160 94.050 ;
        RECT 48.990 89.400 49.160 94.050 ;
        RECT 49.990 89.400 50.160 94.050 ;
        RECT 50.990 89.400 51.160 94.050 ;
        RECT 51.990 89.400 52.160 94.050 ;
        RECT 52.990 89.400 53.160 94.050 ;
        RECT 53.890 89.400 54.060 94.050 ;
        RECT 54.570 89.400 54.740 94.050 ;
        RECT 55.470 89.400 55.640 94.050 ;
        RECT 56.470 89.400 56.640 94.050 ;
        RECT 57.470 89.400 57.640 94.050 ;
        RECT 58.470 89.400 58.640 94.050 ;
        RECT 59.470 89.400 59.640 94.050 ;
        RECT 60.470 89.400 60.640 94.050 ;
        RECT 61.470 89.400 61.640 94.050 ;
        RECT 62.470 89.400 62.640 94.050 ;
        RECT 63.470 89.400 63.640 94.050 ;
        RECT 64.370 89.400 64.540 94.050 ;
        RECT 65.050 89.400 65.220 94.050 ;
        RECT 65.950 89.400 66.120 94.050 ;
        RECT 66.950 89.400 67.120 94.050 ;
        RECT 67.950 89.400 68.120 94.050 ;
        RECT 68.950 89.400 69.120 94.050 ;
        RECT 69.950 89.400 70.120 94.050 ;
        RECT 70.950 89.400 71.120 94.050 ;
        RECT 71.950 89.400 72.120 94.050 ;
        RECT 72.950 89.400 73.120 94.050 ;
        RECT 73.950 89.400 74.120 94.050 ;
        RECT 74.850 89.400 75.020 94.050 ;
        RECT 75.530 89.400 75.700 94.050 ;
        RECT 76.430 89.400 76.600 94.050 ;
        RECT 77.430 89.400 77.600 94.050 ;
        RECT 78.430 89.400 78.600 94.050 ;
        RECT 79.430 89.400 79.600 94.050 ;
        RECT 80.430 89.400 80.600 94.050 ;
        RECT 81.430 89.400 81.600 94.050 ;
        RECT 82.430 89.400 82.600 94.050 ;
        RECT 83.430 89.400 83.600 94.050 ;
        RECT 84.430 89.400 84.600 94.050 ;
        RECT 85.330 89.400 85.500 94.050 ;
        RECT 86.010 89.400 86.180 94.050 ;
        RECT 86.910 89.400 87.080 94.050 ;
        RECT 87.910 89.400 88.080 94.050 ;
        RECT 88.910 89.400 89.080 94.050 ;
        RECT 89.910 89.400 90.080 94.050 ;
        RECT 90.910 89.400 91.080 94.050 ;
        RECT 91.910 89.400 92.080 94.050 ;
        RECT 92.910 89.400 93.080 94.050 ;
        RECT 93.910 89.400 94.080 94.050 ;
        RECT 94.910 89.400 95.080 94.050 ;
        RECT 95.810 89.400 95.980 94.050 ;
        RECT 96.490 89.400 96.660 94.050 ;
        RECT 97.390 89.400 97.560 94.050 ;
        RECT 98.390 89.400 98.560 94.050 ;
        RECT 99.390 89.400 99.560 94.050 ;
        RECT 100.390 89.400 100.560 94.050 ;
        RECT 101.390 89.400 101.560 94.050 ;
        RECT 102.390 89.400 102.560 94.050 ;
        RECT 103.390 89.400 103.560 94.050 ;
        RECT 104.390 89.400 104.560 94.050 ;
        RECT 105.390 89.400 105.560 94.050 ;
        RECT 106.290 89.400 106.460 94.050 ;
        RECT 106.970 89.400 107.140 94.050 ;
        RECT 107.870 89.400 108.040 94.050 ;
        RECT 108.870 89.400 109.040 94.050 ;
        RECT 109.870 89.400 110.040 94.050 ;
        RECT 110.870 89.400 111.040 94.050 ;
        RECT 111.870 89.400 112.040 94.050 ;
        RECT 112.870 89.400 113.040 94.050 ;
        RECT 113.870 89.400 114.040 94.050 ;
        RECT 114.870 89.400 115.040 94.050 ;
        RECT 115.870 89.400 116.040 94.050 ;
        RECT 116.770 89.400 116.940 94.050 ;
        RECT 117.450 88.750 117.750 101.120 ;
        RECT 11.830 88.450 117.750 88.750 ;
        RECT 11.830 87.770 117.750 88.070 ;
        RECT 11.830 75.400 12.130 87.770 ;
        RECT 12.640 82.470 12.810 87.120 ;
        RECT 13.540 82.470 13.710 87.120 ;
        RECT 14.540 82.470 14.710 87.120 ;
        RECT 15.540 82.470 15.710 87.120 ;
        RECT 16.540 82.470 16.710 87.120 ;
        RECT 17.540 82.470 17.710 87.120 ;
        RECT 18.540 82.470 18.710 87.120 ;
        RECT 19.540 82.470 19.710 87.120 ;
        RECT 20.540 82.470 20.710 87.120 ;
        RECT 21.540 82.470 21.710 87.120 ;
        RECT 22.440 82.470 22.610 87.120 ;
        RECT 23.120 82.470 23.290 87.120 ;
        RECT 24.020 82.470 24.190 87.120 ;
        RECT 25.020 82.470 25.190 87.120 ;
        RECT 26.020 82.470 26.190 87.120 ;
        RECT 27.020 82.470 27.190 87.120 ;
        RECT 28.020 82.470 28.190 87.120 ;
        RECT 29.020 82.470 29.190 87.120 ;
        RECT 30.020 82.470 30.190 87.120 ;
        RECT 31.020 82.470 31.190 87.120 ;
        RECT 32.020 82.470 32.190 87.120 ;
        RECT 32.920 82.470 33.090 87.120 ;
        RECT 33.600 82.470 33.770 87.120 ;
        RECT 34.500 82.470 34.670 87.120 ;
        RECT 35.500 82.470 35.670 87.120 ;
        RECT 36.500 82.470 36.670 87.120 ;
        RECT 37.500 82.470 37.670 87.120 ;
        RECT 38.500 82.470 38.670 87.120 ;
        RECT 39.500 82.470 39.670 87.120 ;
        RECT 40.500 82.470 40.670 87.120 ;
        RECT 41.500 82.470 41.670 87.120 ;
        RECT 42.500 82.470 42.670 87.120 ;
        RECT 43.400 82.470 43.570 87.120 ;
        RECT 44.080 82.470 44.250 87.120 ;
        RECT 44.980 82.470 45.150 87.120 ;
        RECT 45.980 82.470 46.150 87.120 ;
        RECT 46.980 82.470 47.150 87.120 ;
        RECT 47.980 82.470 48.150 87.120 ;
        RECT 48.980 82.470 49.150 87.120 ;
        RECT 49.980 82.470 50.150 87.120 ;
        RECT 50.980 82.470 51.150 87.120 ;
        RECT 51.980 82.470 52.150 87.120 ;
        RECT 52.980 82.470 53.150 87.120 ;
        RECT 53.880 82.470 54.050 87.120 ;
        RECT 54.560 82.470 54.730 87.120 ;
        RECT 55.460 82.470 55.630 87.120 ;
        RECT 56.460 82.470 56.630 87.120 ;
        RECT 57.460 82.470 57.630 87.120 ;
        RECT 58.460 82.470 58.630 87.120 ;
        RECT 59.460 82.470 59.630 87.120 ;
        RECT 60.460 82.470 60.630 87.120 ;
        RECT 61.460 82.470 61.630 87.120 ;
        RECT 62.460 82.470 62.630 87.120 ;
        RECT 63.460 82.470 63.630 87.120 ;
        RECT 64.360 82.470 64.530 87.120 ;
        RECT 65.040 82.470 65.210 87.120 ;
        RECT 65.940 82.470 66.110 87.120 ;
        RECT 66.940 82.470 67.110 87.120 ;
        RECT 67.940 82.470 68.110 87.120 ;
        RECT 68.940 82.470 69.110 87.120 ;
        RECT 69.940 82.470 70.110 87.120 ;
        RECT 70.940 82.470 71.110 87.120 ;
        RECT 71.940 82.470 72.110 87.120 ;
        RECT 72.940 82.470 73.110 87.120 ;
        RECT 73.940 82.470 74.110 87.120 ;
        RECT 74.840 82.470 75.010 87.120 ;
        RECT 75.520 82.470 75.690 87.120 ;
        RECT 76.420 82.470 76.590 87.120 ;
        RECT 77.420 82.470 77.590 87.120 ;
        RECT 78.420 82.470 78.590 87.120 ;
        RECT 79.420 82.470 79.590 87.120 ;
        RECT 80.420 82.470 80.590 87.120 ;
        RECT 81.420 82.470 81.590 87.120 ;
        RECT 82.420 82.470 82.590 87.120 ;
        RECT 83.420 82.470 83.590 87.120 ;
        RECT 84.420 82.470 84.590 87.120 ;
        RECT 85.320 82.470 85.490 87.120 ;
        RECT 86.000 82.470 86.170 87.120 ;
        RECT 86.900 82.470 87.070 87.120 ;
        RECT 87.900 82.470 88.070 87.120 ;
        RECT 88.900 82.470 89.070 87.120 ;
        RECT 89.900 82.470 90.070 87.120 ;
        RECT 90.900 82.470 91.070 87.120 ;
        RECT 91.900 82.470 92.070 87.120 ;
        RECT 92.900 82.470 93.070 87.120 ;
        RECT 93.900 82.470 94.070 87.120 ;
        RECT 94.900 82.470 95.070 87.120 ;
        RECT 95.800 82.470 95.970 87.120 ;
        RECT 96.480 82.470 96.650 87.120 ;
        RECT 97.380 82.470 97.550 87.120 ;
        RECT 98.380 82.470 98.550 87.120 ;
        RECT 99.380 82.470 99.550 87.120 ;
        RECT 100.380 82.470 100.550 87.120 ;
        RECT 101.380 82.470 101.550 87.120 ;
        RECT 102.380 82.470 102.550 87.120 ;
        RECT 103.380 82.470 103.550 87.120 ;
        RECT 104.380 82.470 104.550 87.120 ;
        RECT 105.380 82.470 105.550 87.120 ;
        RECT 106.280 82.470 106.450 87.120 ;
        RECT 106.960 82.470 107.130 87.120 ;
        RECT 107.860 82.470 108.030 87.120 ;
        RECT 108.860 82.470 109.030 87.120 ;
        RECT 109.860 82.470 110.030 87.120 ;
        RECT 110.860 82.470 111.030 87.120 ;
        RECT 111.860 82.470 112.030 87.120 ;
        RECT 112.860 82.470 113.030 87.120 ;
        RECT 113.860 82.470 114.030 87.120 ;
        RECT 114.860 82.470 115.030 87.120 ;
        RECT 115.860 82.470 116.030 87.120 ;
        RECT 116.760 82.470 116.930 87.120 ;
        RECT 12.960 81.840 13.290 82.010 ;
        RECT 13.960 81.840 14.290 82.010 ;
        RECT 14.960 81.840 15.290 82.010 ;
        RECT 15.960 81.840 16.290 82.010 ;
        RECT 16.960 81.840 17.290 82.010 ;
        RECT 17.960 81.840 18.290 82.010 ;
        RECT 18.960 81.840 19.290 82.010 ;
        RECT 19.960 81.840 20.290 82.010 ;
        RECT 20.960 81.840 21.290 82.010 ;
        RECT 21.960 81.840 22.290 82.010 ;
        RECT 23.440 81.840 23.770 82.010 ;
        RECT 24.440 81.840 24.770 82.010 ;
        RECT 25.440 81.840 25.770 82.010 ;
        RECT 26.440 81.840 26.770 82.010 ;
        RECT 27.440 81.840 27.770 82.010 ;
        RECT 28.440 81.840 28.770 82.010 ;
        RECT 29.440 81.840 29.770 82.010 ;
        RECT 30.440 81.840 30.770 82.010 ;
        RECT 31.440 81.840 31.770 82.010 ;
        RECT 32.440 81.840 32.770 82.010 ;
        RECT 33.920 81.840 34.250 82.010 ;
        RECT 34.920 81.840 35.250 82.010 ;
        RECT 35.920 81.840 36.250 82.010 ;
        RECT 36.920 81.840 37.250 82.010 ;
        RECT 37.920 81.840 38.250 82.010 ;
        RECT 38.920 81.840 39.250 82.010 ;
        RECT 39.920 81.840 40.250 82.010 ;
        RECT 40.920 81.840 41.250 82.010 ;
        RECT 41.920 81.840 42.250 82.010 ;
        RECT 42.920 81.840 43.250 82.010 ;
        RECT 44.400 81.840 44.730 82.010 ;
        RECT 45.400 81.840 45.730 82.010 ;
        RECT 46.400 81.840 46.730 82.010 ;
        RECT 47.400 81.840 47.730 82.010 ;
        RECT 48.400 81.840 48.730 82.010 ;
        RECT 49.400 81.840 49.730 82.010 ;
        RECT 50.400 81.840 50.730 82.010 ;
        RECT 51.400 81.840 51.730 82.010 ;
        RECT 52.400 81.840 52.730 82.010 ;
        RECT 53.400 81.840 53.730 82.010 ;
        RECT 54.880 81.840 55.210 82.010 ;
        RECT 55.880 81.840 56.210 82.010 ;
        RECT 56.880 81.840 57.210 82.010 ;
        RECT 57.880 81.840 58.210 82.010 ;
        RECT 58.880 81.840 59.210 82.010 ;
        RECT 59.880 81.840 60.210 82.010 ;
        RECT 60.880 81.840 61.210 82.010 ;
        RECT 61.880 81.840 62.210 82.010 ;
        RECT 62.880 81.840 63.210 82.010 ;
        RECT 63.880 81.840 64.210 82.010 ;
        RECT 65.360 81.840 65.690 82.010 ;
        RECT 66.360 81.840 66.690 82.010 ;
        RECT 67.360 81.840 67.690 82.010 ;
        RECT 68.360 81.840 68.690 82.010 ;
        RECT 69.360 81.840 69.690 82.010 ;
        RECT 70.360 81.840 70.690 82.010 ;
        RECT 71.360 81.840 71.690 82.010 ;
        RECT 72.360 81.840 72.690 82.010 ;
        RECT 73.360 81.840 73.690 82.010 ;
        RECT 74.360 81.840 74.690 82.010 ;
        RECT 75.840 81.840 76.170 82.010 ;
        RECT 76.840 81.840 77.170 82.010 ;
        RECT 77.840 81.840 78.170 82.010 ;
        RECT 78.840 81.840 79.170 82.010 ;
        RECT 79.840 81.840 80.170 82.010 ;
        RECT 80.840 81.840 81.170 82.010 ;
        RECT 81.840 81.840 82.170 82.010 ;
        RECT 82.840 81.840 83.170 82.010 ;
        RECT 83.840 81.840 84.170 82.010 ;
        RECT 84.840 81.840 85.170 82.010 ;
        RECT 86.320 81.840 86.650 82.010 ;
        RECT 87.320 81.840 87.650 82.010 ;
        RECT 88.320 81.840 88.650 82.010 ;
        RECT 89.320 81.840 89.650 82.010 ;
        RECT 90.320 81.840 90.650 82.010 ;
        RECT 91.320 81.840 91.650 82.010 ;
        RECT 92.320 81.840 92.650 82.010 ;
        RECT 93.320 81.840 93.650 82.010 ;
        RECT 94.320 81.840 94.650 82.010 ;
        RECT 95.320 81.840 95.650 82.010 ;
        RECT 96.800 81.840 97.130 82.010 ;
        RECT 97.800 81.840 98.130 82.010 ;
        RECT 98.800 81.840 99.130 82.010 ;
        RECT 99.800 81.840 100.130 82.010 ;
        RECT 100.800 81.840 101.130 82.010 ;
        RECT 101.800 81.840 102.130 82.010 ;
        RECT 102.800 81.840 103.130 82.010 ;
        RECT 103.800 81.840 104.130 82.010 ;
        RECT 104.800 81.840 105.130 82.010 ;
        RECT 105.800 81.840 106.130 82.010 ;
        RECT 107.280 81.840 107.610 82.010 ;
        RECT 108.280 81.840 108.610 82.010 ;
        RECT 109.280 81.840 109.610 82.010 ;
        RECT 110.280 81.840 110.610 82.010 ;
        RECT 111.280 81.840 111.610 82.010 ;
        RECT 112.280 81.840 112.610 82.010 ;
        RECT 113.280 81.840 113.610 82.010 ;
        RECT 114.280 81.840 114.610 82.010 ;
        RECT 115.280 81.840 115.610 82.010 ;
        RECT 116.280 81.840 116.610 82.010 ;
        RECT 12.970 81.160 13.300 81.330 ;
        RECT 13.970 81.160 14.300 81.330 ;
        RECT 14.970 81.160 15.300 81.330 ;
        RECT 15.970 81.160 16.300 81.330 ;
        RECT 16.970 81.160 17.300 81.330 ;
        RECT 17.970 81.160 18.300 81.330 ;
        RECT 18.970 81.160 19.300 81.330 ;
        RECT 19.970 81.160 20.300 81.330 ;
        RECT 20.970 81.160 21.300 81.330 ;
        RECT 21.970 81.160 22.300 81.330 ;
        RECT 23.450 81.160 23.780 81.330 ;
        RECT 24.450 81.160 24.780 81.330 ;
        RECT 25.450 81.160 25.780 81.330 ;
        RECT 26.450 81.160 26.780 81.330 ;
        RECT 27.450 81.160 27.780 81.330 ;
        RECT 28.450 81.160 28.780 81.330 ;
        RECT 29.450 81.160 29.780 81.330 ;
        RECT 30.450 81.160 30.780 81.330 ;
        RECT 31.450 81.160 31.780 81.330 ;
        RECT 32.450 81.160 32.780 81.330 ;
        RECT 33.930 81.160 34.260 81.330 ;
        RECT 34.930 81.160 35.260 81.330 ;
        RECT 35.930 81.160 36.260 81.330 ;
        RECT 36.930 81.160 37.260 81.330 ;
        RECT 37.930 81.160 38.260 81.330 ;
        RECT 38.930 81.160 39.260 81.330 ;
        RECT 39.930 81.160 40.260 81.330 ;
        RECT 40.930 81.160 41.260 81.330 ;
        RECT 41.930 81.160 42.260 81.330 ;
        RECT 42.930 81.160 43.260 81.330 ;
        RECT 44.410 81.160 44.740 81.330 ;
        RECT 45.410 81.160 45.740 81.330 ;
        RECT 46.410 81.160 46.740 81.330 ;
        RECT 47.410 81.160 47.740 81.330 ;
        RECT 48.410 81.160 48.740 81.330 ;
        RECT 49.410 81.160 49.740 81.330 ;
        RECT 50.410 81.160 50.740 81.330 ;
        RECT 51.410 81.160 51.740 81.330 ;
        RECT 52.410 81.160 52.740 81.330 ;
        RECT 53.410 81.160 53.740 81.330 ;
        RECT 54.890 81.160 55.220 81.330 ;
        RECT 55.890 81.160 56.220 81.330 ;
        RECT 56.890 81.160 57.220 81.330 ;
        RECT 57.890 81.160 58.220 81.330 ;
        RECT 58.890 81.160 59.220 81.330 ;
        RECT 59.890 81.160 60.220 81.330 ;
        RECT 60.890 81.160 61.220 81.330 ;
        RECT 61.890 81.160 62.220 81.330 ;
        RECT 62.890 81.160 63.220 81.330 ;
        RECT 63.890 81.160 64.220 81.330 ;
        RECT 65.370 81.160 65.700 81.330 ;
        RECT 66.370 81.160 66.700 81.330 ;
        RECT 67.370 81.160 67.700 81.330 ;
        RECT 68.370 81.160 68.700 81.330 ;
        RECT 69.370 81.160 69.700 81.330 ;
        RECT 70.370 81.160 70.700 81.330 ;
        RECT 71.370 81.160 71.700 81.330 ;
        RECT 72.370 81.160 72.700 81.330 ;
        RECT 73.370 81.160 73.700 81.330 ;
        RECT 74.370 81.160 74.700 81.330 ;
        RECT 75.850 81.160 76.180 81.330 ;
        RECT 76.850 81.160 77.180 81.330 ;
        RECT 77.850 81.160 78.180 81.330 ;
        RECT 78.850 81.160 79.180 81.330 ;
        RECT 79.850 81.160 80.180 81.330 ;
        RECT 80.850 81.160 81.180 81.330 ;
        RECT 81.850 81.160 82.180 81.330 ;
        RECT 82.850 81.160 83.180 81.330 ;
        RECT 83.850 81.160 84.180 81.330 ;
        RECT 84.850 81.160 85.180 81.330 ;
        RECT 86.330 81.160 86.660 81.330 ;
        RECT 87.330 81.160 87.660 81.330 ;
        RECT 88.330 81.160 88.660 81.330 ;
        RECT 89.330 81.160 89.660 81.330 ;
        RECT 90.330 81.160 90.660 81.330 ;
        RECT 91.330 81.160 91.660 81.330 ;
        RECT 92.330 81.160 92.660 81.330 ;
        RECT 93.330 81.160 93.660 81.330 ;
        RECT 94.330 81.160 94.660 81.330 ;
        RECT 95.330 81.160 95.660 81.330 ;
        RECT 96.810 81.160 97.140 81.330 ;
        RECT 97.810 81.160 98.140 81.330 ;
        RECT 98.810 81.160 99.140 81.330 ;
        RECT 99.810 81.160 100.140 81.330 ;
        RECT 100.810 81.160 101.140 81.330 ;
        RECT 101.810 81.160 102.140 81.330 ;
        RECT 102.810 81.160 103.140 81.330 ;
        RECT 103.810 81.160 104.140 81.330 ;
        RECT 104.810 81.160 105.140 81.330 ;
        RECT 105.810 81.160 106.140 81.330 ;
        RECT 107.290 81.160 107.620 81.330 ;
        RECT 108.290 81.160 108.620 81.330 ;
        RECT 109.290 81.160 109.620 81.330 ;
        RECT 110.290 81.160 110.620 81.330 ;
        RECT 111.290 81.160 111.620 81.330 ;
        RECT 112.290 81.160 112.620 81.330 ;
        RECT 113.290 81.160 113.620 81.330 ;
        RECT 114.290 81.160 114.620 81.330 ;
        RECT 115.290 81.160 115.620 81.330 ;
        RECT 116.290 81.160 116.620 81.330 ;
        RECT 12.650 76.050 12.820 80.700 ;
        RECT 13.550 76.050 13.720 80.700 ;
        RECT 14.550 76.050 14.720 80.700 ;
        RECT 15.550 76.050 15.720 80.700 ;
        RECT 16.550 76.050 16.720 80.700 ;
        RECT 17.550 76.050 17.720 80.700 ;
        RECT 18.550 76.050 18.720 80.700 ;
        RECT 19.550 76.050 19.720 80.700 ;
        RECT 20.550 76.050 20.720 80.700 ;
        RECT 21.550 76.050 21.720 80.700 ;
        RECT 22.450 76.050 22.620 80.700 ;
        RECT 23.130 76.050 23.300 80.700 ;
        RECT 24.030 76.050 24.200 80.700 ;
        RECT 25.030 76.050 25.200 80.700 ;
        RECT 26.030 76.050 26.200 80.700 ;
        RECT 27.030 76.050 27.200 80.700 ;
        RECT 28.030 76.050 28.200 80.700 ;
        RECT 29.030 76.050 29.200 80.700 ;
        RECT 30.030 76.050 30.200 80.700 ;
        RECT 31.030 76.050 31.200 80.700 ;
        RECT 32.030 76.050 32.200 80.700 ;
        RECT 32.930 76.050 33.100 80.700 ;
        RECT 33.610 76.050 33.780 80.700 ;
        RECT 34.510 76.050 34.680 80.700 ;
        RECT 35.510 76.050 35.680 80.700 ;
        RECT 36.510 76.050 36.680 80.700 ;
        RECT 37.510 76.050 37.680 80.700 ;
        RECT 38.510 76.050 38.680 80.700 ;
        RECT 39.510 76.050 39.680 80.700 ;
        RECT 40.510 76.050 40.680 80.700 ;
        RECT 41.510 76.050 41.680 80.700 ;
        RECT 42.510 76.050 42.680 80.700 ;
        RECT 43.410 76.050 43.580 80.700 ;
        RECT 44.090 76.050 44.260 80.700 ;
        RECT 44.990 76.050 45.160 80.700 ;
        RECT 45.990 76.050 46.160 80.700 ;
        RECT 46.990 76.050 47.160 80.700 ;
        RECT 47.990 76.050 48.160 80.700 ;
        RECT 48.990 76.050 49.160 80.700 ;
        RECT 49.990 76.050 50.160 80.700 ;
        RECT 50.990 76.050 51.160 80.700 ;
        RECT 51.990 76.050 52.160 80.700 ;
        RECT 52.990 76.050 53.160 80.700 ;
        RECT 53.890 76.050 54.060 80.700 ;
        RECT 54.570 76.050 54.740 80.700 ;
        RECT 55.470 76.050 55.640 80.700 ;
        RECT 56.470 76.050 56.640 80.700 ;
        RECT 57.470 76.050 57.640 80.700 ;
        RECT 58.470 76.050 58.640 80.700 ;
        RECT 59.470 76.050 59.640 80.700 ;
        RECT 60.470 76.050 60.640 80.700 ;
        RECT 61.470 76.050 61.640 80.700 ;
        RECT 62.470 76.050 62.640 80.700 ;
        RECT 63.470 76.050 63.640 80.700 ;
        RECT 64.370 76.050 64.540 80.700 ;
        RECT 65.050 76.050 65.220 80.700 ;
        RECT 65.950 76.050 66.120 80.700 ;
        RECT 66.950 76.050 67.120 80.700 ;
        RECT 67.950 76.050 68.120 80.700 ;
        RECT 68.950 76.050 69.120 80.700 ;
        RECT 69.950 76.050 70.120 80.700 ;
        RECT 70.950 76.050 71.120 80.700 ;
        RECT 71.950 76.050 72.120 80.700 ;
        RECT 72.950 76.050 73.120 80.700 ;
        RECT 73.950 76.050 74.120 80.700 ;
        RECT 74.850 76.050 75.020 80.700 ;
        RECT 75.530 76.050 75.700 80.700 ;
        RECT 76.430 76.050 76.600 80.700 ;
        RECT 77.430 76.050 77.600 80.700 ;
        RECT 78.430 76.050 78.600 80.700 ;
        RECT 79.430 76.050 79.600 80.700 ;
        RECT 80.430 76.050 80.600 80.700 ;
        RECT 81.430 76.050 81.600 80.700 ;
        RECT 82.430 76.050 82.600 80.700 ;
        RECT 83.430 76.050 83.600 80.700 ;
        RECT 84.430 76.050 84.600 80.700 ;
        RECT 85.330 76.050 85.500 80.700 ;
        RECT 86.010 76.050 86.180 80.700 ;
        RECT 86.910 76.050 87.080 80.700 ;
        RECT 87.910 76.050 88.080 80.700 ;
        RECT 88.910 76.050 89.080 80.700 ;
        RECT 89.910 76.050 90.080 80.700 ;
        RECT 90.910 76.050 91.080 80.700 ;
        RECT 91.910 76.050 92.080 80.700 ;
        RECT 92.910 76.050 93.080 80.700 ;
        RECT 93.910 76.050 94.080 80.700 ;
        RECT 94.910 76.050 95.080 80.700 ;
        RECT 95.810 76.050 95.980 80.700 ;
        RECT 96.490 76.050 96.660 80.700 ;
        RECT 97.390 76.050 97.560 80.700 ;
        RECT 98.390 76.050 98.560 80.700 ;
        RECT 99.390 76.050 99.560 80.700 ;
        RECT 100.390 76.050 100.560 80.700 ;
        RECT 101.390 76.050 101.560 80.700 ;
        RECT 102.390 76.050 102.560 80.700 ;
        RECT 103.390 76.050 103.560 80.700 ;
        RECT 104.390 76.050 104.560 80.700 ;
        RECT 105.390 76.050 105.560 80.700 ;
        RECT 106.290 76.050 106.460 80.700 ;
        RECT 106.970 76.050 107.140 80.700 ;
        RECT 107.870 76.050 108.040 80.700 ;
        RECT 108.870 76.050 109.040 80.700 ;
        RECT 109.870 76.050 110.040 80.700 ;
        RECT 110.870 76.050 111.040 80.700 ;
        RECT 111.870 76.050 112.040 80.700 ;
        RECT 112.870 76.050 113.040 80.700 ;
        RECT 113.870 76.050 114.040 80.700 ;
        RECT 114.870 76.050 115.040 80.700 ;
        RECT 115.870 76.050 116.040 80.700 ;
        RECT 116.770 76.050 116.940 80.700 ;
        RECT 117.450 75.400 117.750 87.770 ;
        RECT 11.830 75.100 117.750 75.400 ;
        RECT 11.830 74.420 117.750 74.720 ;
        RECT 11.830 62.050 12.130 74.420 ;
        RECT 12.640 69.120 12.810 73.770 ;
        RECT 13.540 69.120 13.710 73.770 ;
        RECT 14.540 69.120 14.710 73.770 ;
        RECT 15.540 69.120 15.710 73.770 ;
        RECT 16.540 69.120 16.710 73.770 ;
        RECT 17.540 69.120 17.710 73.770 ;
        RECT 18.540 69.120 18.710 73.770 ;
        RECT 19.540 69.120 19.710 73.770 ;
        RECT 20.540 69.120 20.710 73.770 ;
        RECT 21.540 69.120 21.710 73.770 ;
        RECT 22.440 69.120 22.610 73.770 ;
        RECT 23.120 69.120 23.290 73.770 ;
        RECT 24.020 69.120 24.190 73.770 ;
        RECT 25.020 69.120 25.190 73.770 ;
        RECT 26.020 69.120 26.190 73.770 ;
        RECT 27.020 69.120 27.190 73.770 ;
        RECT 28.020 69.120 28.190 73.770 ;
        RECT 29.020 69.120 29.190 73.770 ;
        RECT 30.020 69.120 30.190 73.770 ;
        RECT 31.020 69.120 31.190 73.770 ;
        RECT 32.020 69.120 32.190 73.770 ;
        RECT 32.920 69.120 33.090 73.770 ;
        RECT 33.600 69.120 33.770 73.770 ;
        RECT 34.500 69.120 34.670 73.770 ;
        RECT 35.500 69.120 35.670 73.770 ;
        RECT 36.500 69.120 36.670 73.770 ;
        RECT 37.500 69.120 37.670 73.770 ;
        RECT 38.500 69.120 38.670 73.770 ;
        RECT 39.500 69.120 39.670 73.770 ;
        RECT 40.500 69.120 40.670 73.770 ;
        RECT 41.500 69.120 41.670 73.770 ;
        RECT 42.500 69.120 42.670 73.770 ;
        RECT 43.400 69.120 43.570 73.770 ;
        RECT 44.080 69.120 44.250 73.770 ;
        RECT 44.980 69.120 45.150 73.770 ;
        RECT 45.980 69.120 46.150 73.770 ;
        RECT 46.980 69.120 47.150 73.770 ;
        RECT 47.980 69.120 48.150 73.770 ;
        RECT 48.980 69.120 49.150 73.770 ;
        RECT 49.980 69.120 50.150 73.770 ;
        RECT 50.980 69.120 51.150 73.770 ;
        RECT 51.980 69.120 52.150 73.770 ;
        RECT 52.980 69.120 53.150 73.770 ;
        RECT 53.880 69.120 54.050 73.770 ;
        RECT 54.560 69.120 54.730 73.770 ;
        RECT 55.460 69.120 55.630 73.770 ;
        RECT 56.460 69.120 56.630 73.770 ;
        RECT 57.460 69.120 57.630 73.770 ;
        RECT 58.460 69.120 58.630 73.770 ;
        RECT 59.460 69.120 59.630 73.770 ;
        RECT 60.460 69.120 60.630 73.770 ;
        RECT 61.460 69.120 61.630 73.770 ;
        RECT 62.460 69.120 62.630 73.770 ;
        RECT 63.460 69.120 63.630 73.770 ;
        RECT 64.360 69.120 64.530 73.770 ;
        RECT 65.040 69.120 65.210 73.770 ;
        RECT 65.940 69.120 66.110 73.770 ;
        RECT 66.940 69.120 67.110 73.770 ;
        RECT 67.940 69.120 68.110 73.770 ;
        RECT 68.940 69.120 69.110 73.770 ;
        RECT 69.940 69.120 70.110 73.770 ;
        RECT 70.940 69.120 71.110 73.770 ;
        RECT 71.940 69.120 72.110 73.770 ;
        RECT 72.940 69.120 73.110 73.770 ;
        RECT 73.940 69.120 74.110 73.770 ;
        RECT 74.840 69.120 75.010 73.770 ;
        RECT 75.520 69.120 75.690 73.770 ;
        RECT 76.420 69.120 76.590 73.770 ;
        RECT 77.420 69.120 77.590 73.770 ;
        RECT 78.420 69.120 78.590 73.770 ;
        RECT 79.420 69.120 79.590 73.770 ;
        RECT 80.420 69.120 80.590 73.770 ;
        RECT 81.420 69.120 81.590 73.770 ;
        RECT 82.420 69.120 82.590 73.770 ;
        RECT 83.420 69.120 83.590 73.770 ;
        RECT 84.420 69.120 84.590 73.770 ;
        RECT 85.320 69.120 85.490 73.770 ;
        RECT 86.000 69.120 86.170 73.770 ;
        RECT 86.900 69.120 87.070 73.770 ;
        RECT 87.900 69.120 88.070 73.770 ;
        RECT 88.900 69.120 89.070 73.770 ;
        RECT 89.900 69.120 90.070 73.770 ;
        RECT 90.900 69.120 91.070 73.770 ;
        RECT 91.900 69.120 92.070 73.770 ;
        RECT 92.900 69.120 93.070 73.770 ;
        RECT 93.900 69.120 94.070 73.770 ;
        RECT 94.900 69.120 95.070 73.770 ;
        RECT 95.800 69.120 95.970 73.770 ;
        RECT 96.480 69.120 96.650 73.770 ;
        RECT 97.380 69.120 97.550 73.770 ;
        RECT 98.380 69.120 98.550 73.770 ;
        RECT 99.380 69.120 99.550 73.770 ;
        RECT 100.380 69.120 100.550 73.770 ;
        RECT 101.380 69.120 101.550 73.770 ;
        RECT 102.380 69.120 102.550 73.770 ;
        RECT 103.380 69.120 103.550 73.770 ;
        RECT 104.380 69.120 104.550 73.770 ;
        RECT 105.380 69.120 105.550 73.770 ;
        RECT 106.280 69.120 106.450 73.770 ;
        RECT 106.960 69.120 107.130 73.770 ;
        RECT 107.860 69.120 108.030 73.770 ;
        RECT 108.860 69.120 109.030 73.770 ;
        RECT 109.860 69.120 110.030 73.770 ;
        RECT 110.860 69.120 111.030 73.770 ;
        RECT 111.860 69.120 112.030 73.770 ;
        RECT 112.860 69.120 113.030 73.770 ;
        RECT 113.860 69.120 114.030 73.770 ;
        RECT 114.860 69.120 115.030 73.770 ;
        RECT 115.860 69.120 116.030 73.770 ;
        RECT 116.760 69.120 116.930 73.770 ;
        RECT 12.960 68.490 13.290 68.660 ;
        RECT 13.960 68.490 14.290 68.660 ;
        RECT 14.960 68.490 15.290 68.660 ;
        RECT 15.960 68.490 16.290 68.660 ;
        RECT 16.960 68.490 17.290 68.660 ;
        RECT 17.960 68.490 18.290 68.660 ;
        RECT 18.960 68.490 19.290 68.660 ;
        RECT 19.960 68.490 20.290 68.660 ;
        RECT 20.960 68.490 21.290 68.660 ;
        RECT 21.960 68.490 22.290 68.660 ;
        RECT 23.440 68.490 23.770 68.660 ;
        RECT 24.440 68.490 24.770 68.660 ;
        RECT 25.440 68.490 25.770 68.660 ;
        RECT 26.440 68.490 26.770 68.660 ;
        RECT 27.440 68.490 27.770 68.660 ;
        RECT 28.440 68.490 28.770 68.660 ;
        RECT 29.440 68.490 29.770 68.660 ;
        RECT 30.440 68.490 30.770 68.660 ;
        RECT 31.440 68.490 31.770 68.660 ;
        RECT 32.440 68.490 32.770 68.660 ;
        RECT 33.920 68.490 34.250 68.660 ;
        RECT 34.920 68.490 35.250 68.660 ;
        RECT 35.920 68.490 36.250 68.660 ;
        RECT 36.920 68.490 37.250 68.660 ;
        RECT 37.920 68.490 38.250 68.660 ;
        RECT 38.920 68.490 39.250 68.660 ;
        RECT 39.920 68.490 40.250 68.660 ;
        RECT 40.920 68.490 41.250 68.660 ;
        RECT 41.920 68.490 42.250 68.660 ;
        RECT 42.920 68.490 43.250 68.660 ;
        RECT 44.400 68.490 44.730 68.660 ;
        RECT 45.400 68.490 45.730 68.660 ;
        RECT 46.400 68.490 46.730 68.660 ;
        RECT 47.400 68.490 47.730 68.660 ;
        RECT 48.400 68.490 48.730 68.660 ;
        RECT 49.400 68.490 49.730 68.660 ;
        RECT 50.400 68.490 50.730 68.660 ;
        RECT 51.400 68.490 51.730 68.660 ;
        RECT 52.400 68.490 52.730 68.660 ;
        RECT 53.400 68.490 53.730 68.660 ;
        RECT 54.880 68.490 55.210 68.660 ;
        RECT 55.880 68.490 56.210 68.660 ;
        RECT 56.880 68.490 57.210 68.660 ;
        RECT 57.880 68.490 58.210 68.660 ;
        RECT 58.880 68.490 59.210 68.660 ;
        RECT 59.880 68.490 60.210 68.660 ;
        RECT 60.880 68.490 61.210 68.660 ;
        RECT 61.880 68.490 62.210 68.660 ;
        RECT 62.880 68.490 63.210 68.660 ;
        RECT 63.880 68.490 64.210 68.660 ;
        RECT 65.360 68.490 65.690 68.660 ;
        RECT 66.360 68.490 66.690 68.660 ;
        RECT 67.360 68.490 67.690 68.660 ;
        RECT 68.360 68.490 68.690 68.660 ;
        RECT 69.360 68.490 69.690 68.660 ;
        RECT 70.360 68.490 70.690 68.660 ;
        RECT 71.360 68.490 71.690 68.660 ;
        RECT 72.360 68.490 72.690 68.660 ;
        RECT 73.360 68.490 73.690 68.660 ;
        RECT 74.360 68.490 74.690 68.660 ;
        RECT 75.840 68.490 76.170 68.660 ;
        RECT 76.840 68.490 77.170 68.660 ;
        RECT 77.840 68.490 78.170 68.660 ;
        RECT 78.840 68.490 79.170 68.660 ;
        RECT 79.840 68.490 80.170 68.660 ;
        RECT 80.840 68.490 81.170 68.660 ;
        RECT 81.840 68.490 82.170 68.660 ;
        RECT 82.840 68.490 83.170 68.660 ;
        RECT 83.840 68.490 84.170 68.660 ;
        RECT 84.840 68.490 85.170 68.660 ;
        RECT 86.320 68.490 86.650 68.660 ;
        RECT 87.320 68.490 87.650 68.660 ;
        RECT 88.320 68.490 88.650 68.660 ;
        RECT 89.320 68.490 89.650 68.660 ;
        RECT 90.320 68.490 90.650 68.660 ;
        RECT 91.320 68.490 91.650 68.660 ;
        RECT 92.320 68.490 92.650 68.660 ;
        RECT 93.320 68.490 93.650 68.660 ;
        RECT 94.320 68.490 94.650 68.660 ;
        RECT 95.320 68.490 95.650 68.660 ;
        RECT 96.800 68.490 97.130 68.660 ;
        RECT 97.800 68.490 98.130 68.660 ;
        RECT 98.800 68.490 99.130 68.660 ;
        RECT 99.800 68.490 100.130 68.660 ;
        RECT 100.800 68.490 101.130 68.660 ;
        RECT 101.800 68.490 102.130 68.660 ;
        RECT 102.800 68.490 103.130 68.660 ;
        RECT 103.800 68.490 104.130 68.660 ;
        RECT 104.800 68.490 105.130 68.660 ;
        RECT 105.800 68.490 106.130 68.660 ;
        RECT 107.280 68.490 107.610 68.660 ;
        RECT 108.280 68.490 108.610 68.660 ;
        RECT 109.280 68.490 109.610 68.660 ;
        RECT 110.280 68.490 110.610 68.660 ;
        RECT 111.280 68.490 111.610 68.660 ;
        RECT 112.280 68.490 112.610 68.660 ;
        RECT 113.280 68.490 113.610 68.660 ;
        RECT 114.280 68.490 114.610 68.660 ;
        RECT 115.280 68.490 115.610 68.660 ;
        RECT 116.280 68.490 116.610 68.660 ;
        RECT 12.970 67.810 13.300 67.980 ;
        RECT 13.970 67.810 14.300 67.980 ;
        RECT 14.970 67.810 15.300 67.980 ;
        RECT 15.970 67.810 16.300 67.980 ;
        RECT 16.970 67.810 17.300 67.980 ;
        RECT 17.970 67.810 18.300 67.980 ;
        RECT 18.970 67.810 19.300 67.980 ;
        RECT 19.970 67.810 20.300 67.980 ;
        RECT 20.970 67.810 21.300 67.980 ;
        RECT 21.970 67.810 22.300 67.980 ;
        RECT 23.450 67.810 23.780 67.980 ;
        RECT 24.450 67.810 24.780 67.980 ;
        RECT 25.450 67.810 25.780 67.980 ;
        RECT 26.450 67.810 26.780 67.980 ;
        RECT 27.450 67.810 27.780 67.980 ;
        RECT 28.450 67.810 28.780 67.980 ;
        RECT 29.450 67.810 29.780 67.980 ;
        RECT 30.450 67.810 30.780 67.980 ;
        RECT 31.450 67.810 31.780 67.980 ;
        RECT 32.450 67.810 32.780 67.980 ;
        RECT 33.930 67.810 34.260 67.980 ;
        RECT 34.930 67.810 35.260 67.980 ;
        RECT 35.930 67.810 36.260 67.980 ;
        RECT 36.930 67.810 37.260 67.980 ;
        RECT 37.930 67.810 38.260 67.980 ;
        RECT 38.930 67.810 39.260 67.980 ;
        RECT 39.930 67.810 40.260 67.980 ;
        RECT 40.930 67.810 41.260 67.980 ;
        RECT 41.930 67.810 42.260 67.980 ;
        RECT 42.930 67.810 43.260 67.980 ;
        RECT 44.410 67.810 44.740 67.980 ;
        RECT 45.410 67.810 45.740 67.980 ;
        RECT 46.410 67.810 46.740 67.980 ;
        RECT 47.410 67.810 47.740 67.980 ;
        RECT 48.410 67.810 48.740 67.980 ;
        RECT 49.410 67.810 49.740 67.980 ;
        RECT 50.410 67.810 50.740 67.980 ;
        RECT 51.410 67.810 51.740 67.980 ;
        RECT 52.410 67.810 52.740 67.980 ;
        RECT 53.410 67.810 53.740 67.980 ;
        RECT 54.890 67.810 55.220 67.980 ;
        RECT 55.890 67.810 56.220 67.980 ;
        RECT 56.890 67.810 57.220 67.980 ;
        RECT 57.890 67.810 58.220 67.980 ;
        RECT 58.890 67.810 59.220 67.980 ;
        RECT 59.890 67.810 60.220 67.980 ;
        RECT 60.890 67.810 61.220 67.980 ;
        RECT 61.890 67.810 62.220 67.980 ;
        RECT 62.890 67.810 63.220 67.980 ;
        RECT 63.890 67.810 64.220 67.980 ;
        RECT 65.370 67.810 65.700 67.980 ;
        RECT 66.370 67.810 66.700 67.980 ;
        RECT 67.370 67.810 67.700 67.980 ;
        RECT 68.370 67.810 68.700 67.980 ;
        RECT 69.370 67.810 69.700 67.980 ;
        RECT 70.370 67.810 70.700 67.980 ;
        RECT 71.370 67.810 71.700 67.980 ;
        RECT 72.370 67.810 72.700 67.980 ;
        RECT 73.370 67.810 73.700 67.980 ;
        RECT 74.370 67.810 74.700 67.980 ;
        RECT 75.850 67.810 76.180 67.980 ;
        RECT 76.850 67.810 77.180 67.980 ;
        RECT 77.850 67.810 78.180 67.980 ;
        RECT 78.850 67.810 79.180 67.980 ;
        RECT 79.850 67.810 80.180 67.980 ;
        RECT 80.850 67.810 81.180 67.980 ;
        RECT 81.850 67.810 82.180 67.980 ;
        RECT 82.850 67.810 83.180 67.980 ;
        RECT 83.850 67.810 84.180 67.980 ;
        RECT 84.850 67.810 85.180 67.980 ;
        RECT 86.330 67.810 86.660 67.980 ;
        RECT 87.330 67.810 87.660 67.980 ;
        RECT 88.330 67.810 88.660 67.980 ;
        RECT 89.330 67.810 89.660 67.980 ;
        RECT 90.330 67.810 90.660 67.980 ;
        RECT 91.330 67.810 91.660 67.980 ;
        RECT 92.330 67.810 92.660 67.980 ;
        RECT 93.330 67.810 93.660 67.980 ;
        RECT 94.330 67.810 94.660 67.980 ;
        RECT 95.330 67.810 95.660 67.980 ;
        RECT 96.810 67.810 97.140 67.980 ;
        RECT 97.810 67.810 98.140 67.980 ;
        RECT 98.810 67.810 99.140 67.980 ;
        RECT 99.810 67.810 100.140 67.980 ;
        RECT 100.810 67.810 101.140 67.980 ;
        RECT 101.810 67.810 102.140 67.980 ;
        RECT 102.810 67.810 103.140 67.980 ;
        RECT 103.810 67.810 104.140 67.980 ;
        RECT 104.810 67.810 105.140 67.980 ;
        RECT 105.810 67.810 106.140 67.980 ;
        RECT 107.290 67.810 107.620 67.980 ;
        RECT 108.290 67.810 108.620 67.980 ;
        RECT 109.290 67.810 109.620 67.980 ;
        RECT 110.290 67.810 110.620 67.980 ;
        RECT 111.290 67.810 111.620 67.980 ;
        RECT 112.290 67.810 112.620 67.980 ;
        RECT 113.290 67.810 113.620 67.980 ;
        RECT 114.290 67.810 114.620 67.980 ;
        RECT 115.290 67.810 115.620 67.980 ;
        RECT 116.290 67.810 116.620 67.980 ;
        RECT 12.650 62.700 12.820 67.350 ;
        RECT 13.550 62.700 13.720 67.350 ;
        RECT 14.550 62.700 14.720 67.350 ;
        RECT 15.550 62.700 15.720 67.350 ;
        RECT 16.550 62.700 16.720 67.350 ;
        RECT 17.550 62.700 17.720 67.350 ;
        RECT 18.550 62.700 18.720 67.350 ;
        RECT 19.550 62.700 19.720 67.350 ;
        RECT 20.550 62.700 20.720 67.350 ;
        RECT 21.550 62.700 21.720 67.350 ;
        RECT 22.450 62.700 22.620 67.350 ;
        RECT 23.130 62.700 23.300 67.350 ;
        RECT 24.030 62.700 24.200 67.350 ;
        RECT 25.030 62.700 25.200 67.350 ;
        RECT 26.030 62.700 26.200 67.350 ;
        RECT 27.030 62.700 27.200 67.350 ;
        RECT 28.030 62.700 28.200 67.350 ;
        RECT 29.030 62.700 29.200 67.350 ;
        RECT 30.030 62.700 30.200 67.350 ;
        RECT 31.030 62.700 31.200 67.350 ;
        RECT 32.030 62.700 32.200 67.350 ;
        RECT 32.930 62.700 33.100 67.350 ;
        RECT 33.610 62.700 33.780 67.350 ;
        RECT 34.510 62.700 34.680 67.350 ;
        RECT 35.510 62.700 35.680 67.350 ;
        RECT 36.510 62.700 36.680 67.350 ;
        RECT 37.510 62.700 37.680 67.350 ;
        RECT 38.510 62.700 38.680 67.350 ;
        RECT 39.510 62.700 39.680 67.350 ;
        RECT 40.510 62.700 40.680 67.350 ;
        RECT 41.510 62.700 41.680 67.350 ;
        RECT 42.510 62.700 42.680 67.350 ;
        RECT 43.410 62.700 43.580 67.350 ;
        RECT 44.090 62.700 44.260 67.350 ;
        RECT 44.990 62.700 45.160 67.350 ;
        RECT 45.990 62.700 46.160 67.350 ;
        RECT 46.990 62.700 47.160 67.350 ;
        RECT 47.990 62.700 48.160 67.350 ;
        RECT 48.990 62.700 49.160 67.350 ;
        RECT 49.990 62.700 50.160 67.350 ;
        RECT 50.990 62.700 51.160 67.350 ;
        RECT 51.990 62.700 52.160 67.350 ;
        RECT 52.990 62.700 53.160 67.350 ;
        RECT 53.890 62.700 54.060 67.350 ;
        RECT 54.570 62.700 54.740 67.350 ;
        RECT 55.470 62.700 55.640 67.350 ;
        RECT 56.470 62.700 56.640 67.350 ;
        RECT 57.470 62.700 57.640 67.350 ;
        RECT 58.470 62.700 58.640 67.350 ;
        RECT 59.470 62.700 59.640 67.350 ;
        RECT 60.470 62.700 60.640 67.350 ;
        RECT 61.470 62.700 61.640 67.350 ;
        RECT 62.470 62.700 62.640 67.350 ;
        RECT 63.470 62.700 63.640 67.350 ;
        RECT 64.370 62.700 64.540 67.350 ;
        RECT 65.050 62.700 65.220 67.350 ;
        RECT 65.950 62.700 66.120 67.350 ;
        RECT 66.950 62.700 67.120 67.350 ;
        RECT 67.950 62.700 68.120 67.350 ;
        RECT 68.950 62.700 69.120 67.350 ;
        RECT 69.950 62.700 70.120 67.350 ;
        RECT 70.950 62.700 71.120 67.350 ;
        RECT 71.950 62.700 72.120 67.350 ;
        RECT 72.950 62.700 73.120 67.350 ;
        RECT 73.950 62.700 74.120 67.350 ;
        RECT 74.850 62.700 75.020 67.350 ;
        RECT 75.530 62.700 75.700 67.350 ;
        RECT 76.430 62.700 76.600 67.350 ;
        RECT 77.430 62.700 77.600 67.350 ;
        RECT 78.430 62.700 78.600 67.350 ;
        RECT 79.430 62.700 79.600 67.350 ;
        RECT 80.430 62.700 80.600 67.350 ;
        RECT 81.430 62.700 81.600 67.350 ;
        RECT 82.430 62.700 82.600 67.350 ;
        RECT 83.430 62.700 83.600 67.350 ;
        RECT 84.430 62.700 84.600 67.350 ;
        RECT 85.330 62.700 85.500 67.350 ;
        RECT 86.010 62.700 86.180 67.350 ;
        RECT 86.910 62.700 87.080 67.350 ;
        RECT 87.910 62.700 88.080 67.350 ;
        RECT 88.910 62.700 89.080 67.350 ;
        RECT 89.910 62.700 90.080 67.350 ;
        RECT 90.910 62.700 91.080 67.350 ;
        RECT 91.910 62.700 92.080 67.350 ;
        RECT 92.910 62.700 93.080 67.350 ;
        RECT 93.910 62.700 94.080 67.350 ;
        RECT 94.910 62.700 95.080 67.350 ;
        RECT 95.810 62.700 95.980 67.350 ;
        RECT 96.490 62.700 96.660 67.350 ;
        RECT 97.390 62.700 97.560 67.350 ;
        RECT 98.390 62.700 98.560 67.350 ;
        RECT 99.390 62.700 99.560 67.350 ;
        RECT 100.390 62.700 100.560 67.350 ;
        RECT 101.390 62.700 101.560 67.350 ;
        RECT 102.390 62.700 102.560 67.350 ;
        RECT 103.390 62.700 103.560 67.350 ;
        RECT 104.390 62.700 104.560 67.350 ;
        RECT 105.390 62.700 105.560 67.350 ;
        RECT 106.290 62.700 106.460 67.350 ;
        RECT 106.970 62.700 107.140 67.350 ;
        RECT 107.870 62.700 108.040 67.350 ;
        RECT 108.870 62.700 109.040 67.350 ;
        RECT 109.870 62.700 110.040 67.350 ;
        RECT 110.870 62.700 111.040 67.350 ;
        RECT 111.870 62.700 112.040 67.350 ;
        RECT 112.870 62.700 113.040 67.350 ;
        RECT 113.870 62.700 114.040 67.350 ;
        RECT 114.870 62.700 115.040 67.350 ;
        RECT 115.870 62.700 116.040 67.350 ;
        RECT 116.770 62.700 116.940 67.350 ;
        RECT 117.450 62.050 117.750 74.420 ;
        RECT 11.830 61.750 117.750 62.050 ;
        RECT 52.130 11.580 63.730 11.880 ;
        RECT 52.130 5.300 52.430 11.580 ;
        RECT 53.270 11.060 53.600 11.230 ;
        RECT 54.270 11.060 54.600 11.230 ;
        RECT 55.270 11.060 55.600 11.230 ;
        RECT 56.270 11.060 56.600 11.230 ;
        RECT 57.270 11.060 57.600 11.230 ;
        RECT 58.270 11.060 58.600 11.230 ;
        RECT 59.270 11.060 59.600 11.230 ;
        RECT 60.270 11.060 60.600 11.230 ;
        RECT 61.270 11.060 61.600 11.230 ;
        RECT 62.270 11.060 62.600 11.230 ;
        RECT 52.950 5.950 53.120 10.600 ;
        RECT 53.850 5.950 54.020 10.600 ;
        RECT 54.850 5.950 55.020 10.600 ;
        RECT 55.850 5.950 56.020 10.600 ;
        RECT 56.850 5.950 57.020 10.600 ;
        RECT 57.850 5.950 58.020 10.600 ;
        RECT 58.850 5.950 59.020 10.600 ;
        RECT 59.850 5.950 60.020 10.600 ;
        RECT 60.850 5.950 61.020 10.600 ;
        RECT 61.850 5.950 62.020 10.600 ;
        RECT 62.750 5.950 62.920 10.600 ;
        RECT 63.430 5.300 63.730 11.580 ;
        RECT 52.130 5.000 63.730 5.300 ;
        RECT 64.020 11.580 75.620 11.880 ;
        RECT 64.020 5.300 64.320 11.580 ;
        RECT 65.160 11.060 65.490 11.230 ;
        RECT 66.160 11.060 66.490 11.230 ;
        RECT 67.160 11.060 67.490 11.230 ;
        RECT 68.160 11.060 68.490 11.230 ;
        RECT 69.160 11.060 69.490 11.230 ;
        RECT 70.160 11.060 70.490 11.230 ;
        RECT 71.160 11.060 71.490 11.230 ;
        RECT 72.160 11.060 72.490 11.230 ;
        RECT 73.160 11.060 73.490 11.230 ;
        RECT 74.160 11.060 74.490 11.230 ;
        RECT 64.840 5.950 65.010 10.600 ;
        RECT 65.740 5.950 65.910 10.600 ;
        RECT 66.740 5.950 66.910 10.600 ;
        RECT 67.740 5.950 67.910 10.600 ;
        RECT 68.740 5.950 68.910 10.600 ;
        RECT 69.740 5.950 69.910 10.600 ;
        RECT 70.740 5.950 70.910 10.600 ;
        RECT 71.740 5.950 71.910 10.600 ;
        RECT 72.740 5.950 72.910 10.600 ;
        RECT 73.740 5.950 73.910 10.600 ;
        RECT 74.640 5.950 74.810 10.600 ;
        RECT 75.320 5.300 75.620 11.580 ;
        RECT 64.020 5.000 75.620 5.300 ;
      LAYER met1 ;
        RECT 4.000 11.880 6.000 220.760 ;
        RECT 118.980 172.480 142.440 172.710 ;
        RECT 118.980 119.480 119.210 172.480 ;
        RECT 120.850 171.200 140.580 171.900 ;
        RECT 119.660 121.190 120.460 170.800 ;
        RECT 140.970 121.190 141.770 170.800 ;
        RECT 120.850 120.100 140.580 120.800 ;
        RECT 142.210 119.480 142.440 172.480 ;
        RECT 118.980 119.250 142.440 119.480 ;
        RECT 11.830 114.470 117.750 114.770 ;
        RECT 11.830 102.100 12.130 114.470 ;
        RECT 12.560 109.190 12.880 113.800 ;
        RECT 13.510 109.190 13.740 114.470 ;
        RECT 14.460 109.190 14.780 113.800 ;
        RECT 15.510 109.190 15.740 114.470 ;
        RECT 16.460 109.190 16.780 113.800 ;
        RECT 17.510 109.190 17.740 114.470 ;
        RECT 18.460 109.190 18.780 113.800 ;
        RECT 19.510 109.190 19.740 114.470 ;
        RECT 20.460 109.190 20.780 113.800 ;
        RECT 21.510 109.190 21.740 114.470 ;
        RECT 22.410 109.190 23.320 113.800 ;
        RECT 23.990 109.190 24.220 114.470 ;
        RECT 24.940 109.190 25.260 113.800 ;
        RECT 25.990 109.190 26.220 114.470 ;
        RECT 26.940 109.190 27.260 113.800 ;
        RECT 27.990 109.190 28.220 114.470 ;
        RECT 28.940 109.190 29.260 113.800 ;
        RECT 29.990 109.190 30.220 114.470 ;
        RECT 30.940 109.190 31.260 113.800 ;
        RECT 31.990 109.190 32.220 114.470 ;
        RECT 32.890 109.190 33.800 113.800 ;
        RECT 34.470 109.190 34.700 114.470 ;
        RECT 35.420 109.190 35.740 113.800 ;
        RECT 36.470 109.190 36.700 114.470 ;
        RECT 37.420 109.190 37.740 113.800 ;
        RECT 38.470 109.190 38.700 114.470 ;
        RECT 39.420 109.190 39.740 113.800 ;
        RECT 40.470 109.190 40.700 114.470 ;
        RECT 41.420 109.190 41.740 113.800 ;
        RECT 42.470 109.190 42.700 114.470 ;
        RECT 43.370 109.190 44.280 113.800 ;
        RECT 44.950 109.190 45.180 114.470 ;
        RECT 45.900 109.190 46.220 113.800 ;
        RECT 46.950 109.190 47.180 114.470 ;
        RECT 47.900 109.190 48.220 113.800 ;
        RECT 48.950 109.190 49.180 114.470 ;
        RECT 49.900 109.190 50.220 113.800 ;
        RECT 50.950 109.190 51.180 114.470 ;
        RECT 51.900 109.190 52.220 113.800 ;
        RECT 52.950 109.190 53.180 114.470 ;
        RECT 53.850 109.190 54.760 113.800 ;
        RECT 55.430 109.190 55.660 114.470 ;
        RECT 56.380 109.190 56.700 113.800 ;
        RECT 57.430 109.190 57.660 114.470 ;
        RECT 58.380 109.190 58.700 113.800 ;
        RECT 59.430 109.190 59.660 114.470 ;
        RECT 60.380 109.190 60.700 113.800 ;
        RECT 61.430 109.190 61.660 114.470 ;
        RECT 62.380 109.190 62.700 113.800 ;
        RECT 63.430 109.190 63.660 114.470 ;
        RECT 64.330 109.190 65.240 113.800 ;
        RECT 65.910 109.190 66.140 114.470 ;
        RECT 66.860 109.190 67.180 113.800 ;
        RECT 67.910 109.190 68.140 114.470 ;
        RECT 68.860 109.190 69.180 113.800 ;
        RECT 69.910 109.190 70.140 114.470 ;
        RECT 70.860 109.190 71.180 113.800 ;
        RECT 71.910 109.190 72.140 114.470 ;
        RECT 72.860 109.190 73.180 113.800 ;
        RECT 73.910 109.190 74.140 114.470 ;
        RECT 74.810 109.190 75.720 113.800 ;
        RECT 76.390 109.190 76.620 114.470 ;
        RECT 77.340 109.190 77.660 113.800 ;
        RECT 78.390 109.190 78.620 114.470 ;
        RECT 79.340 109.190 79.660 113.800 ;
        RECT 80.390 109.190 80.620 114.470 ;
        RECT 81.340 109.190 81.660 113.800 ;
        RECT 82.390 109.190 82.620 114.470 ;
        RECT 83.340 109.190 83.660 113.800 ;
        RECT 84.390 109.190 84.620 114.470 ;
        RECT 85.290 109.190 86.200 113.800 ;
        RECT 86.870 109.190 87.100 114.470 ;
        RECT 87.820 109.190 88.140 113.800 ;
        RECT 88.870 109.190 89.100 114.470 ;
        RECT 89.820 109.190 90.140 113.800 ;
        RECT 90.870 109.190 91.100 114.470 ;
        RECT 91.820 109.190 92.140 113.800 ;
        RECT 92.870 109.190 93.100 114.470 ;
        RECT 93.820 109.190 94.140 113.800 ;
        RECT 94.870 109.190 95.100 114.470 ;
        RECT 95.770 109.190 96.680 113.800 ;
        RECT 97.350 109.190 97.580 114.470 ;
        RECT 98.300 109.190 98.620 113.800 ;
        RECT 99.350 109.190 99.580 114.470 ;
        RECT 100.300 109.190 100.620 113.800 ;
        RECT 101.350 109.190 101.580 114.470 ;
        RECT 102.300 109.190 102.620 113.800 ;
        RECT 103.350 109.190 103.580 114.470 ;
        RECT 104.300 109.190 104.620 113.800 ;
        RECT 105.350 109.190 105.580 114.470 ;
        RECT 106.250 109.190 107.160 113.800 ;
        RECT 107.830 109.190 108.060 114.470 ;
        RECT 108.780 109.190 109.100 113.800 ;
        RECT 109.830 109.190 110.060 114.470 ;
        RECT 110.780 109.190 111.100 113.800 ;
        RECT 111.830 109.190 112.060 114.470 ;
        RECT 112.780 109.190 113.100 113.800 ;
        RECT 113.830 109.190 114.060 114.470 ;
        RECT 114.780 109.190 115.100 113.800 ;
        RECT 115.830 109.190 116.060 114.470 ;
        RECT 116.730 109.190 117.050 113.800 ;
        RECT 12.950 107.830 116.630 108.740 ;
        RECT 12.570 102.770 12.890 107.380 ;
        RECT 13.520 102.100 13.750 107.380 ;
        RECT 14.470 102.770 14.790 107.380 ;
        RECT 15.520 102.100 15.750 107.380 ;
        RECT 16.470 102.770 16.790 107.380 ;
        RECT 17.520 102.100 17.750 107.380 ;
        RECT 18.470 102.770 18.790 107.380 ;
        RECT 19.520 102.100 19.750 107.380 ;
        RECT 20.470 102.770 20.790 107.380 ;
        RECT 21.520 102.100 21.750 107.380 ;
        RECT 22.420 102.770 23.330 107.380 ;
        RECT 24.000 102.100 24.230 107.380 ;
        RECT 24.950 102.770 25.270 107.380 ;
        RECT 26.000 102.100 26.230 107.380 ;
        RECT 26.950 102.770 27.270 107.380 ;
        RECT 28.000 102.100 28.230 107.380 ;
        RECT 28.950 102.770 29.270 107.380 ;
        RECT 30.000 102.100 30.230 107.380 ;
        RECT 30.950 102.770 31.270 107.380 ;
        RECT 32.000 102.100 32.230 107.380 ;
        RECT 32.900 102.770 33.810 107.380 ;
        RECT 34.480 102.100 34.710 107.380 ;
        RECT 35.430 102.770 35.750 107.380 ;
        RECT 36.480 102.100 36.710 107.380 ;
        RECT 37.430 102.770 37.750 107.380 ;
        RECT 38.480 102.100 38.710 107.380 ;
        RECT 39.430 102.770 39.750 107.380 ;
        RECT 40.480 102.100 40.710 107.380 ;
        RECT 41.430 102.770 41.750 107.380 ;
        RECT 42.480 102.100 42.710 107.380 ;
        RECT 43.380 102.770 44.290 107.380 ;
        RECT 44.960 102.100 45.190 107.380 ;
        RECT 45.910 102.770 46.230 107.380 ;
        RECT 46.960 102.100 47.190 107.380 ;
        RECT 47.910 102.770 48.230 107.380 ;
        RECT 48.960 102.100 49.190 107.380 ;
        RECT 49.910 102.770 50.230 107.380 ;
        RECT 50.960 102.100 51.190 107.380 ;
        RECT 51.910 102.770 52.230 107.380 ;
        RECT 52.960 102.100 53.190 107.380 ;
        RECT 53.860 102.770 54.770 107.380 ;
        RECT 55.440 102.100 55.670 107.380 ;
        RECT 56.390 102.770 56.710 107.380 ;
        RECT 57.440 102.100 57.670 107.380 ;
        RECT 58.390 102.770 58.710 107.380 ;
        RECT 59.440 102.100 59.670 107.380 ;
        RECT 60.390 102.770 60.710 107.380 ;
        RECT 61.440 102.100 61.670 107.380 ;
        RECT 62.390 102.770 62.710 107.380 ;
        RECT 63.440 102.100 63.670 107.380 ;
        RECT 64.340 102.770 65.250 107.380 ;
        RECT 65.920 102.100 66.150 107.380 ;
        RECT 66.870 102.770 67.190 107.380 ;
        RECT 67.920 102.100 68.150 107.380 ;
        RECT 68.870 102.770 69.190 107.380 ;
        RECT 69.920 102.100 70.150 107.380 ;
        RECT 70.870 102.770 71.190 107.380 ;
        RECT 71.920 102.100 72.150 107.380 ;
        RECT 72.870 102.770 73.190 107.380 ;
        RECT 73.920 102.100 74.150 107.380 ;
        RECT 74.820 102.770 75.730 107.380 ;
        RECT 76.400 102.100 76.630 107.380 ;
        RECT 77.350 102.770 77.670 107.380 ;
        RECT 78.400 102.100 78.630 107.380 ;
        RECT 79.350 102.770 79.670 107.380 ;
        RECT 80.400 102.100 80.630 107.380 ;
        RECT 81.350 102.770 81.670 107.380 ;
        RECT 82.400 102.100 82.630 107.380 ;
        RECT 83.350 102.770 83.670 107.380 ;
        RECT 84.400 102.100 84.630 107.380 ;
        RECT 85.300 102.770 86.210 107.380 ;
        RECT 86.880 102.100 87.110 107.380 ;
        RECT 87.830 102.770 88.150 107.380 ;
        RECT 88.880 102.100 89.110 107.380 ;
        RECT 89.830 102.770 90.150 107.380 ;
        RECT 90.880 102.100 91.110 107.380 ;
        RECT 91.830 102.770 92.150 107.380 ;
        RECT 92.880 102.100 93.110 107.380 ;
        RECT 93.830 102.770 94.150 107.380 ;
        RECT 94.880 102.100 95.110 107.380 ;
        RECT 95.780 102.770 96.690 107.380 ;
        RECT 97.360 102.100 97.590 107.380 ;
        RECT 98.310 102.770 98.630 107.380 ;
        RECT 99.360 102.100 99.590 107.380 ;
        RECT 100.310 102.770 100.630 107.380 ;
        RECT 101.360 102.100 101.590 107.380 ;
        RECT 102.310 102.770 102.630 107.380 ;
        RECT 103.360 102.100 103.590 107.380 ;
        RECT 104.310 102.770 104.630 107.380 ;
        RECT 105.360 102.100 105.590 107.380 ;
        RECT 106.260 102.770 107.170 107.380 ;
        RECT 107.840 102.100 108.070 107.380 ;
        RECT 108.790 102.770 109.110 107.380 ;
        RECT 109.840 102.100 110.070 107.380 ;
        RECT 110.790 102.770 111.110 107.380 ;
        RECT 111.840 102.100 112.070 107.380 ;
        RECT 112.790 102.770 113.110 107.380 ;
        RECT 113.840 102.100 114.070 107.380 ;
        RECT 114.790 102.770 115.110 107.380 ;
        RECT 115.840 102.100 116.070 107.380 ;
        RECT 116.740 102.780 117.060 107.380 ;
        RECT 116.740 102.770 116.970 102.780 ;
        RECT 117.450 102.100 117.750 114.470 ;
        RECT 11.830 101.120 117.750 102.100 ;
        RECT 11.830 88.750 12.130 101.120 ;
        RECT 12.560 95.840 12.880 100.450 ;
        RECT 13.510 95.840 13.740 101.120 ;
        RECT 14.460 95.840 14.780 100.450 ;
        RECT 15.510 95.840 15.740 101.120 ;
        RECT 16.460 95.840 16.780 100.450 ;
        RECT 17.510 95.840 17.740 101.120 ;
        RECT 18.460 95.840 18.780 100.450 ;
        RECT 19.510 95.840 19.740 101.120 ;
        RECT 20.460 95.840 20.780 100.450 ;
        RECT 21.510 95.840 21.740 101.120 ;
        RECT 22.410 95.840 23.320 100.450 ;
        RECT 23.990 95.840 24.220 101.120 ;
        RECT 24.940 95.840 25.260 100.450 ;
        RECT 25.990 95.840 26.220 101.120 ;
        RECT 26.940 95.840 27.260 100.450 ;
        RECT 27.990 95.840 28.220 101.120 ;
        RECT 28.940 95.840 29.260 100.450 ;
        RECT 29.990 95.840 30.220 101.120 ;
        RECT 30.940 95.840 31.260 100.450 ;
        RECT 31.990 95.840 32.220 101.120 ;
        RECT 32.890 95.840 33.800 100.450 ;
        RECT 34.470 95.840 34.700 101.120 ;
        RECT 35.420 95.840 35.740 100.450 ;
        RECT 36.470 95.840 36.700 101.120 ;
        RECT 37.420 95.840 37.740 100.450 ;
        RECT 38.470 95.840 38.700 101.120 ;
        RECT 39.420 95.840 39.740 100.450 ;
        RECT 40.470 95.840 40.700 101.120 ;
        RECT 41.420 95.840 41.740 100.450 ;
        RECT 42.470 95.840 42.700 101.120 ;
        RECT 43.370 95.840 44.280 100.450 ;
        RECT 44.950 95.840 45.180 101.120 ;
        RECT 45.900 95.840 46.220 100.450 ;
        RECT 46.950 95.840 47.180 101.120 ;
        RECT 47.900 95.840 48.220 100.450 ;
        RECT 48.950 95.840 49.180 101.120 ;
        RECT 49.900 95.840 50.220 100.450 ;
        RECT 50.950 95.840 51.180 101.120 ;
        RECT 51.900 95.840 52.220 100.450 ;
        RECT 52.950 95.840 53.180 101.120 ;
        RECT 53.850 95.840 54.760 100.450 ;
        RECT 55.430 95.840 55.660 101.120 ;
        RECT 56.380 95.840 56.700 100.450 ;
        RECT 57.430 95.840 57.660 101.120 ;
        RECT 58.380 95.840 58.700 100.450 ;
        RECT 59.430 95.840 59.660 101.120 ;
        RECT 60.380 95.840 60.700 100.450 ;
        RECT 61.430 95.840 61.660 101.120 ;
        RECT 62.380 95.840 62.700 100.450 ;
        RECT 63.430 95.840 63.660 101.120 ;
        RECT 64.330 95.840 65.240 100.450 ;
        RECT 65.910 95.840 66.140 101.120 ;
        RECT 66.860 95.840 67.180 100.450 ;
        RECT 67.910 95.840 68.140 101.120 ;
        RECT 68.860 95.840 69.180 100.450 ;
        RECT 69.910 95.840 70.140 101.120 ;
        RECT 70.860 95.840 71.180 100.450 ;
        RECT 71.910 95.840 72.140 101.120 ;
        RECT 72.860 95.840 73.180 100.450 ;
        RECT 73.910 95.840 74.140 101.120 ;
        RECT 74.810 95.840 75.720 100.450 ;
        RECT 76.390 95.840 76.620 101.120 ;
        RECT 77.340 95.840 77.660 100.450 ;
        RECT 78.390 95.840 78.620 101.120 ;
        RECT 79.340 95.840 79.660 100.450 ;
        RECT 80.390 95.840 80.620 101.120 ;
        RECT 81.340 95.840 81.660 100.450 ;
        RECT 82.390 95.840 82.620 101.120 ;
        RECT 83.340 95.840 83.660 100.450 ;
        RECT 84.390 95.840 84.620 101.120 ;
        RECT 85.290 95.840 86.200 100.450 ;
        RECT 86.870 95.840 87.100 101.120 ;
        RECT 87.820 95.840 88.140 100.450 ;
        RECT 88.870 95.840 89.100 101.120 ;
        RECT 89.820 95.840 90.140 100.450 ;
        RECT 90.870 95.840 91.100 101.120 ;
        RECT 91.820 95.840 92.140 100.450 ;
        RECT 92.870 95.840 93.100 101.120 ;
        RECT 93.820 95.840 94.140 100.450 ;
        RECT 94.870 95.840 95.100 101.120 ;
        RECT 95.770 95.840 96.680 100.450 ;
        RECT 97.350 95.840 97.580 101.120 ;
        RECT 98.300 95.840 98.620 100.450 ;
        RECT 99.350 95.840 99.580 101.120 ;
        RECT 100.300 95.840 100.620 100.450 ;
        RECT 101.350 95.840 101.580 101.120 ;
        RECT 102.300 95.840 102.620 100.450 ;
        RECT 103.350 95.840 103.580 101.120 ;
        RECT 104.300 95.840 104.620 100.450 ;
        RECT 105.350 95.840 105.580 101.120 ;
        RECT 106.250 95.840 107.160 100.450 ;
        RECT 107.830 95.840 108.060 101.120 ;
        RECT 108.780 95.840 109.100 100.450 ;
        RECT 109.830 95.840 110.060 101.120 ;
        RECT 110.780 95.840 111.100 100.450 ;
        RECT 111.830 95.840 112.060 101.120 ;
        RECT 112.780 95.840 113.100 100.450 ;
        RECT 113.830 95.840 114.060 101.120 ;
        RECT 114.780 95.840 115.100 100.450 ;
        RECT 115.830 95.840 116.060 101.120 ;
        RECT 116.730 95.840 117.050 100.450 ;
        RECT 12.950 94.480 116.630 95.390 ;
        RECT 12.570 89.420 12.890 94.030 ;
        RECT 13.520 88.750 13.750 94.030 ;
        RECT 14.470 89.420 14.790 94.030 ;
        RECT 15.520 88.750 15.750 94.030 ;
        RECT 16.470 89.420 16.790 94.030 ;
        RECT 17.520 88.750 17.750 94.030 ;
        RECT 18.470 89.420 18.790 94.030 ;
        RECT 19.520 88.750 19.750 94.030 ;
        RECT 20.470 89.420 20.790 94.030 ;
        RECT 21.520 88.750 21.750 94.030 ;
        RECT 22.420 89.420 23.330 94.030 ;
        RECT 24.000 88.750 24.230 94.030 ;
        RECT 24.950 89.420 25.270 94.030 ;
        RECT 26.000 88.750 26.230 94.030 ;
        RECT 26.950 89.420 27.270 94.030 ;
        RECT 28.000 88.750 28.230 94.030 ;
        RECT 28.950 89.420 29.270 94.030 ;
        RECT 30.000 88.750 30.230 94.030 ;
        RECT 30.950 89.420 31.270 94.030 ;
        RECT 32.000 88.750 32.230 94.030 ;
        RECT 32.900 89.420 33.810 94.030 ;
        RECT 34.480 88.750 34.710 94.030 ;
        RECT 35.430 89.420 35.750 94.030 ;
        RECT 36.480 88.750 36.710 94.030 ;
        RECT 37.430 89.420 37.750 94.030 ;
        RECT 38.480 88.750 38.710 94.030 ;
        RECT 39.430 89.420 39.750 94.030 ;
        RECT 40.480 88.750 40.710 94.030 ;
        RECT 41.430 89.420 41.750 94.030 ;
        RECT 42.480 88.750 42.710 94.030 ;
        RECT 43.380 89.420 44.290 94.030 ;
        RECT 44.960 88.750 45.190 94.030 ;
        RECT 45.910 89.420 46.230 94.030 ;
        RECT 46.960 88.750 47.190 94.030 ;
        RECT 47.910 89.420 48.230 94.030 ;
        RECT 48.960 88.750 49.190 94.030 ;
        RECT 49.910 89.420 50.230 94.030 ;
        RECT 50.960 88.750 51.190 94.030 ;
        RECT 51.910 89.420 52.230 94.030 ;
        RECT 52.960 88.750 53.190 94.030 ;
        RECT 53.860 89.420 54.770 94.030 ;
        RECT 55.440 88.750 55.670 94.030 ;
        RECT 56.390 89.420 56.710 94.030 ;
        RECT 57.440 88.750 57.670 94.030 ;
        RECT 58.390 89.420 58.710 94.030 ;
        RECT 59.440 88.750 59.670 94.030 ;
        RECT 60.390 89.420 60.710 94.030 ;
        RECT 61.440 88.750 61.670 94.030 ;
        RECT 62.390 89.420 62.710 94.030 ;
        RECT 63.440 88.750 63.670 94.030 ;
        RECT 64.340 89.420 65.250 94.030 ;
        RECT 65.920 88.750 66.150 94.030 ;
        RECT 66.870 89.420 67.190 94.030 ;
        RECT 67.920 88.750 68.150 94.030 ;
        RECT 68.870 89.420 69.190 94.030 ;
        RECT 69.920 88.750 70.150 94.030 ;
        RECT 70.870 89.420 71.190 94.030 ;
        RECT 71.920 88.750 72.150 94.030 ;
        RECT 72.870 89.420 73.190 94.030 ;
        RECT 73.920 88.750 74.150 94.030 ;
        RECT 74.820 89.420 75.730 94.030 ;
        RECT 76.400 88.750 76.630 94.030 ;
        RECT 77.350 89.420 77.670 94.030 ;
        RECT 78.400 88.750 78.630 94.030 ;
        RECT 79.350 89.420 79.670 94.030 ;
        RECT 80.400 88.750 80.630 94.030 ;
        RECT 81.350 89.420 81.670 94.030 ;
        RECT 82.400 88.750 82.630 94.030 ;
        RECT 83.350 89.420 83.670 94.030 ;
        RECT 84.400 88.750 84.630 94.030 ;
        RECT 85.300 89.420 86.210 94.030 ;
        RECT 86.880 88.750 87.110 94.030 ;
        RECT 87.830 89.420 88.150 94.030 ;
        RECT 88.880 88.750 89.110 94.030 ;
        RECT 89.830 89.420 90.150 94.030 ;
        RECT 90.880 88.750 91.110 94.030 ;
        RECT 91.830 89.420 92.150 94.030 ;
        RECT 92.880 88.750 93.110 94.030 ;
        RECT 93.830 89.420 94.150 94.030 ;
        RECT 94.880 88.750 95.110 94.030 ;
        RECT 95.780 89.420 96.690 94.030 ;
        RECT 97.360 88.750 97.590 94.030 ;
        RECT 98.310 89.420 98.630 94.030 ;
        RECT 99.360 88.750 99.590 94.030 ;
        RECT 100.310 89.420 100.630 94.030 ;
        RECT 101.360 88.750 101.590 94.030 ;
        RECT 102.310 89.420 102.630 94.030 ;
        RECT 103.360 88.750 103.590 94.030 ;
        RECT 104.310 89.420 104.630 94.030 ;
        RECT 105.360 88.750 105.590 94.030 ;
        RECT 106.260 89.420 107.170 94.030 ;
        RECT 107.840 88.750 108.070 94.030 ;
        RECT 108.790 89.420 109.110 94.030 ;
        RECT 109.840 88.750 110.070 94.030 ;
        RECT 110.790 89.420 111.110 94.030 ;
        RECT 111.840 88.750 112.070 94.030 ;
        RECT 112.790 89.420 113.110 94.030 ;
        RECT 113.840 88.750 114.070 94.030 ;
        RECT 114.790 89.420 115.110 94.030 ;
        RECT 115.840 88.750 116.070 94.030 ;
        RECT 116.740 89.430 117.060 94.030 ;
        RECT 116.740 89.420 116.970 89.430 ;
        RECT 117.450 88.750 117.750 101.120 ;
        RECT 11.830 87.770 117.750 88.750 ;
        RECT 11.830 75.400 12.130 87.770 ;
        RECT 12.560 82.490 12.880 87.100 ;
        RECT 13.510 82.490 13.740 87.770 ;
        RECT 14.460 82.490 14.780 87.100 ;
        RECT 15.510 82.490 15.740 87.770 ;
        RECT 16.460 82.490 16.780 87.100 ;
        RECT 17.510 82.490 17.740 87.770 ;
        RECT 18.460 82.490 18.780 87.100 ;
        RECT 19.510 82.490 19.740 87.770 ;
        RECT 20.460 82.490 20.780 87.100 ;
        RECT 21.510 82.490 21.740 87.770 ;
        RECT 22.410 82.490 23.320 87.100 ;
        RECT 23.990 82.490 24.220 87.770 ;
        RECT 24.940 82.490 25.260 87.100 ;
        RECT 25.990 82.490 26.220 87.770 ;
        RECT 26.940 82.490 27.260 87.100 ;
        RECT 27.990 82.490 28.220 87.770 ;
        RECT 28.940 82.490 29.260 87.100 ;
        RECT 29.990 82.490 30.220 87.770 ;
        RECT 30.940 82.490 31.260 87.100 ;
        RECT 31.990 82.490 32.220 87.770 ;
        RECT 32.890 82.490 33.800 87.100 ;
        RECT 34.470 82.490 34.700 87.770 ;
        RECT 35.420 82.490 35.740 87.100 ;
        RECT 36.470 82.490 36.700 87.770 ;
        RECT 37.420 82.490 37.740 87.100 ;
        RECT 38.470 82.490 38.700 87.770 ;
        RECT 39.420 82.490 39.740 87.100 ;
        RECT 40.470 82.490 40.700 87.770 ;
        RECT 41.420 82.490 41.740 87.100 ;
        RECT 42.470 82.490 42.700 87.770 ;
        RECT 43.370 82.490 44.280 87.100 ;
        RECT 44.950 82.490 45.180 87.770 ;
        RECT 45.900 82.490 46.220 87.100 ;
        RECT 46.950 82.490 47.180 87.770 ;
        RECT 47.900 82.490 48.220 87.100 ;
        RECT 48.950 82.490 49.180 87.770 ;
        RECT 49.900 82.490 50.220 87.100 ;
        RECT 50.950 82.490 51.180 87.770 ;
        RECT 51.900 82.490 52.220 87.100 ;
        RECT 52.950 82.490 53.180 87.770 ;
        RECT 53.850 82.490 54.760 87.100 ;
        RECT 55.430 82.490 55.660 87.770 ;
        RECT 56.380 82.490 56.700 87.100 ;
        RECT 57.430 82.490 57.660 87.770 ;
        RECT 58.380 82.490 58.700 87.100 ;
        RECT 59.430 82.490 59.660 87.770 ;
        RECT 60.380 82.490 60.700 87.100 ;
        RECT 61.430 82.490 61.660 87.770 ;
        RECT 62.380 82.490 62.700 87.100 ;
        RECT 63.430 82.490 63.660 87.770 ;
        RECT 64.330 82.490 65.240 87.100 ;
        RECT 65.910 82.490 66.140 87.770 ;
        RECT 66.860 82.490 67.180 87.100 ;
        RECT 67.910 82.490 68.140 87.770 ;
        RECT 68.860 82.490 69.180 87.100 ;
        RECT 69.910 82.490 70.140 87.770 ;
        RECT 70.860 82.490 71.180 87.100 ;
        RECT 71.910 82.490 72.140 87.770 ;
        RECT 72.860 82.490 73.180 87.100 ;
        RECT 73.910 82.490 74.140 87.770 ;
        RECT 74.810 82.490 75.720 87.100 ;
        RECT 76.390 82.490 76.620 87.770 ;
        RECT 77.340 82.490 77.660 87.100 ;
        RECT 78.390 82.490 78.620 87.770 ;
        RECT 79.340 82.490 79.660 87.100 ;
        RECT 80.390 82.490 80.620 87.770 ;
        RECT 81.340 82.490 81.660 87.100 ;
        RECT 82.390 82.490 82.620 87.770 ;
        RECT 83.340 82.490 83.660 87.100 ;
        RECT 84.390 82.490 84.620 87.770 ;
        RECT 85.290 82.490 86.200 87.100 ;
        RECT 86.870 82.490 87.100 87.770 ;
        RECT 87.820 82.490 88.140 87.100 ;
        RECT 88.870 82.490 89.100 87.770 ;
        RECT 89.820 82.490 90.140 87.100 ;
        RECT 90.870 82.490 91.100 87.770 ;
        RECT 91.820 82.490 92.140 87.100 ;
        RECT 92.870 82.490 93.100 87.770 ;
        RECT 93.820 82.490 94.140 87.100 ;
        RECT 94.870 82.490 95.100 87.770 ;
        RECT 95.770 82.490 96.680 87.100 ;
        RECT 97.350 82.490 97.580 87.770 ;
        RECT 98.300 82.490 98.620 87.100 ;
        RECT 99.350 82.490 99.580 87.770 ;
        RECT 100.300 82.490 100.620 87.100 ;
        RECT 101.350 82.490 101.580 87.770 ;
        RECT 102.300 82.490 102.620 87.100 ;
        RECT 103.350 82.490 103.580 87.770 ;
        RECT 104.300 82.490 104.620 87.100 ;
        RECT 105.350 82.490 105.580 87.770 ;
        RECT 106.250 82.490 107.160 87.100 ;
        RECT 107.830 82.490 108.060 87.770 ;
        RECT 108.780 82.490 109.100 87.100 ;
        RECT 109.830 82.490 110.060 87.770 ;
        RECT 110.780 82.490 111.100 87.100 ;
        RECT 111.830 82.490 112.060 87.770 ;
        RECT 112.780 82.490 113.100 87.100 ;
        RECT 113.830 82.490 114.060 87.770 ;
        RECT 114.780 82.490 115.100 87.100 ;
        RECT 115.830 82.490 116.060 87.770 ;
        RECT 116.730 82.490 117.050 87.100 ;
        RECT 12.950 81.130 116.630 82.040 ;
        RECT 12.570 76.070 12.890 80.680 ;
        RECT 13.520 75.400 13.750 80.680 ;
        RECT 14.470 76.070 14.790 80.680 ;
        RECT 15.520 75.400 15.750 80.680 ;
        RECT 16.470 76.070 16.790 80.680 ;
        RECT 17.520 75.400 17.750 80.680 ;
        RECT 18.470 76.070 18.790 80.680 ;
        RECT 19.520 75.400 19.750 80.680 ;
        RECT 20.470 76.070 20.790 80.680 ;
        RECT 21.520 75.400 21.750 80.680 ;
        RECT 22.420 76.070 23.330 80.680 ;
        RECT 24.000 75.400 24.230 80.680 ;
        RECT 24.950 76.070 25.270 80.680 ;
        RECT 26.000 75.400 26.230 80.680 ;
        RECT 26.950 76.070 27.270 80.680 ;
        RECT 28.000 75.400 28.230 80.680 ;
        RECT 28.950 76.070 29.270 80.680 ;
        RECT 30.000 75.400 30.230 80.680 ;
        RECT 30.950 76.070 31.270 80.680 ;
        RECT 32.000 75.400 32.230 80.680 ;
        RECT 32.900 76.070 33.810 80.680 ;
        RECT 34.480 75.400 34.710 80.680 ;
        RECT 35.430 76.070 35.750 80.680 ;
        RECT 36.480 75.400 36.710 80.680 ;
        RECT 37.430 76.070 37.750 80.680 ;
        RECT 38.480 75.400 38.710 80.680 ;
        RECT 39.430 76.070 39.750 80.680 ;
        RECT 40.480 75.400 40.710 80.680 ;
        RECT 41.430 76.070 41.750 80.680 ;
        RECT 42.480 75.400 42.710 80.680 ;
        RECT 43.380 76.070 44.290 80.680 ;
        RECT 44.960 75.400 45.190 80.680 ;
        RECT 45.910 76.070 46.230 80.680 ;
        RECT 46.960 75.400 47.190 80.680 ;
        RECT 47.910 76.070 48.230 80.680 ;
        RECT 48.960 75.400 49.190 80.680 ;
        RECT 49.910 76.070 50.230 80.680 ;
        RECT 50.960 75.400 51.190 80.680 ;
        RECT 51.910 76.070 52.230 80.680 ;
        RECT 52.960 75.400 53.190 80.680 ;
        RECT 53.860 76.070 54.770 80.680 ;
        RECT 55.440 75.400 55.670 80.680 ;
        RECT 56.390 76.070 56.710 80.680 ;
        RECT 57.440 75.400 57.670 80.680 ;
        RECT 58.390 76.070 58.710 80.680 ;
        RECT 59.440 75.400 59.670 80.680 ;
        RECT 60.390 76.070 60.710 80.680 ;
        RECT 61.440 75.400 61.670 80.680 ;
        RECT 62.390 76.070 62.710 80.680 ;
        RECT 63.440 75.400 63.670 80.680 ;
        RECT 64.340 76.070 65.250 80.680 ;
        RECT 65.920 75.400 66.150 80.680 ;
        RECT 66.870 76.070 67.190 80.680 ;
        RECT 67.920 75.400 68.150 80.680 ;
        RECT 68.870 76.070 69.190 80.680 ;
        RECT 69.920 75.400 70.150 80.680 ;
        RECT 70.870 76.070 71.190 80.680 ;
        RECT 71.920 75.400 72.150 80.680 ;
        RECT 72.870 76.070 73.190 80.680 ;
        RECT 73.920 75.400 74.150 80.680 ;
        RECT 74.820 76.070 75.730 80.680 ;
        RECT 76.400 75.400 76.630 80.680 ;
        RECT 77.350 76.070 77.670 80.680 ;
        RECT 78.400 75.400 78.630 80.680 ;
        RECT 79.350 76.070 79.670 80.680 ;
        RECT 80.400 75.400 80.630 80.680 ;
        RECT 81.350 76.070 81.670 80.680 ;
        RECT 82.400 75.400 82.630 80.680 ;
        RECT 83.350 76.070 83.670 80.680 ;
        RECT 84.400 75.400 84.630 80.680 ;
        RECT 85.300 76.070 86.210 80.680 ;
        RECT 86.880 75.400 87.110 80.680 ;
        RECT 87.830 76.070 88.150 80.680 ;
        RECT 88.880 75.400 89.110 80.680 ;
        RECT 89.830 76.070 90.150 80.680 ;
        RECT 90.880 75.400 91.110 80.680 ;
        RECT 91.830 76.070 92.150 80.680 ;
        RECT 92.880 75.400 93.110 80.680 ;
        RECT 93.830 76.070 94.150 80.680 ;
        RECT 94.880 75.400 95.110 80.680 ;
        RECT 95.780 76.070 96.690 80.680 ;
        RECT 97.360 75.400 97.590 80.680 ;
        RECT 98.310 76.070 98.630 80.680 ;
        RECT 99.360 75.400 99.590 80.680 ;
        RECT 100.310 76.070 100.630 80.680 ;
        RECT 101.360 75.400 101.590 80.680 ;
        RECT 102.310 76.070 102.630 80.680 ;
        RECT 103.360 75.400 103.590 80.680 ;
        RECT 104.310 76.070 104.630 80.680 ;
        RECT 105.360 75.400 105.590 80.680 ;
        RECT 106.260 76.070 107.170 80.680 ;
        RECT 107.840 75.400 108.070 80.680 ;
        RECT 108.790 76.070 109.110 80.680 ;
        RECT 109.840 75.400 110.070 80.680 ;
        RECT 110.790 76.070 111.110 80.680 ;
        RECT 111.840 75.400 112.070 80.680 ;
        RECT 112.790 76.070 113.110 80.680 ;
        RECT 113.840 75.400 114.070 80.680 ;
        RECT 114.790 76.070 115.110 80.680 ;
        RECT 115.840 75.400 116.070 80.680 ;
        RECT 116.740 76.080 117.060 80.680 ;
        RECT 116.740 76.070 116.970 76.080 ;
        RECT 117.450 75.400 117.750 87.770 ;
        RECT 11.830 74.420 117.750 75.400 ;
        RECT 11.830 62.050 12.130 74.420 ;
        RECT 12.560 69.140 12.880 73.750 ;
        RECT 13.510 69.140 13.740 74.420 ;
        RECT 14.460 69.140 14.780 73.750 ;
        RECT 15.510 69.140 15.740 74.420 ;
        RECT 16.460 69.140 16.780 73.750 ;
        RECT 17.510 69.140 17.740 74.420 ;
        RECT 18.460 69.140 18.780 73.750 ;
        RECT 19.510 69.140 19.740 74.420 ;
        RECT 20.460 69.140 20.780 73.750 ;
        RECT 21.510 69.140 21.740 74.420 ;
        RECT 22.410 69.140 23.320 73.750 ;
        RECT 23.990 69.140 24.220 74.420 ;
        RECT 24.940 69.140 25.260 73.750 ;
        RECT 25.990 69.140 26.220 74.420 ;
        RECT 26.940 69.140 27.260 73.750 ;
        RECT 27.990 69.140 28.220 74.420 ;
        RECT 28.940 69.140 29.260 73.750 ;
        RECT 29.990 69.140 30.220 74.420 ;
        RECT 30.940 69.140 31.260 73.750 ;
        RECT 31.990 69.140 32.220 74.420 ;
        RECT 32.890 69.140 33.800 73.750 ;
        RECT 34.470 69.140 34.700 74.420 ;
        RECT 35.420 69.140 35.740 73.750 ;
        RECT 36.470 69.140 36.700 74.420 ;
        RECT 37.420 69.140 37.740 73.750 ;
        RECT 38.470 69.140 38.700 74.420 ;
        RECT 39.420 69.140 39.740 73.750 ;
        RECT 40.470 69.140 40.700 74.420 ;
        RECT 41.420 69.140 41.740 73.750 ;
        RECT 42.470 69.140 42.700 74.420 ;
        RECT 43.370 69.140 44.280 73.750 ;
        RECT 44.950 69.140 45.180 74.420 ;
        RECT 45.900 69.140 46.220 73.750 ;
        RECT 46.950 69.140 47.180 74.420 ;
        RECT 47.900 69.140 48.220 73.750 ;
        RECT 48.950 69.140 49.180 74.420 ;
        RECT 49.900 69.140 50.220 73.750 ;
        RECT 50.950 69.140 51.180 74.420 ;
        RECT 51.900 69.140 52.220 73.750 ;
        RECT 52.950 69.140 53.180 74.420 ;
        RECT 53.850 69.140 54.760 73.750 ;
        RECT 55.430 69.140 55.660 74.420 ;
        RECT 56.380 69.140 56.700 73.750 ;
        RECT 57.430 69.140 57.660 74.420 ;
        RECT 58.380 69.140 58.700 73.750 ;
        RECT 59.430 69.140 59.660 74.420 ;
        RECT 60.380 69.140 60.700 73.750 ;
        RECT 61.430 69.140 61.660 74.420 ;
        RECT 62.380 69.140 62.700 73.750 ;
        RECT 63.430 69.140 63.660 74.420 ;
        RECT 64.330 69.140 65.240 73.750 ;
        RECT 65.910 69.140 66.140 74.420 ;
        RECT 66.860 69.140 67.180 73.750 ;
        RECT 67.910 69.140 68.140 74.420 ;
        RECT 68.860 69.140 69.180 73.750 ;
        RECT 69.910 69.140 70.140 74.420 ;
        RECT 70.860 69.140 71.180 73.750 ;
        RECT 71.910 69.140 72.140 74.420 ;
        RECT 72.860 69.140 73.180 73.750 ;
        RECT 73.910 69.140 74.140 74.420 ;
        RECT 74.810 69.140 75.720 73.750 ;
        RECT 76.390 69.140 76.620 74.420 ;
        RECT 77.340 69.140 77.660 73.750 ;
        RECT 78.390 69.140 78.620 74.420 ;
        RECT 79.340 69.140 79.660 73.750 ;
        RECT 80.390 69.140 80.620 74.420 ;
        RECT 81.340 69.140 81.660 73.750 ;
        RECT 82.390 69.140 82.620 74.420 ;
        RECT 83.340 69.140 83.660 73.750 ;
        RECT 84.390 69.140 84.620 74.420 ;
        RECT 85.290 69.140 86.200 73.750 ;
        RECT 86.870 69.140 87.100 74.420 ;
        RECT 87.820 69.140 88.140 73.750 ;
        RECT 88.870 69.140 89.100 74.420 ;
        RECT 89.820 69.140 90.140 73.750 ;
        RECT 90.870 69.140 91.100 74.420 ;
        RECT 91.820 69.140 92.140 73.750 ;
        RECT 92.870 69.140 93.100 74.420 ;
        RECT 93.820 69.140 94.140 73.750 ;
        RECT 94.870 69.140 95.100 74.420 ;
        RECT 95.770 69.140 96.680 73.750 ;
        RECT 97.350 69.140 97.580 74.420 ;
        RECT 98.300 69.140 98.620 73.750 ;
        RECT 99.350 69.140 99.580 74.420 ;
        RECT 100.300 69.140 100.620 73.750 ;
        RECT 101.350 69.140 101.580 74.420 ;
        RECT 102.300 69.140 102.620 73.750 ;
        RECT 103.350 69.140 103.580 74.420 ;
        RECT 104.300 69.140 104.620 73.750 ;
        RECT 105.350 69.140 105.580 74.420 ;
        RECT 106.250 69.140 107.160 73.750 ;
        RECT 107.830 69.140 108.060 74.420 ;
        RECT 108.780 69.140 109.100 73.750 ;
        RECT 109.830 69.140 110.060 74.420 ;
        RECT 110.780 69.140 111.100 73.750 ;
        RECT 111.830 69.140 112.060 74.420 ;
        RECT 112.780 69.140 113.100 73.750 ;
        RECT 113.830 69.140 114.060 74.420 ;
        RECT 114.780 69.140 115.100 73.750 ;
        RECT 115.830 69.140 116.060 74.420 ;
        RECT 116.730 69.140 117.050 73.750 ;
        RECT 12.950 67.780 116.630 68.690 ;
        RECT 12.570 62.720 12.890 67.330 ;
        RECT 13.520 62.050 13.750 67.330 ;
        RECT 14.470 62.720 14.790 67.330 ;
        RECT 15.520 62.050 15.750 67.330 ;
        RECT 16.470 62.720 16.790 67.330 ;
        RECT 17.520 62.050 17.750 67.330 ;
        RECT 18.470 62.720 18.790 67.330 ;
        RECT 19.520 62.050 19.750 67.330 ;
        RECT 20.470 62.720 20.790 67.330 ;
        RECT 21.520 62.050 21.750 67.330 ;
        RECT 22.420 62.720 23.330 67.330 ;
        RECT 24.000 62.050 24.230 67.330 ;
        RECT 24.950 62.720 25.270 67.330 ;
        RECT 26.000 62.050 26.230 67.330 ;
        RECT 26.950 62.720 27.270 67.330 ;
        RECT 28.000 62.050 28.230 67.330 ;
        RECT 28.950 62.720 29.270 67.330 ;
        RECT 30.000 62.050 30.230 67.330 ;
        RECT 30.950 62.720 31.270 67.330 ;
        RECT 32.000 62.050 32.230 67.330 ;
        RECT 32.900 62.720 33.810 67.330 ;
        RECT 34.480 62.050 34.710 67.330 ;
        RECT 35.430 62.720 35.750 67.330 ;
        RECT 36.480 62.050 36.710 67.330 ;
        RECT 37.430 62.720 37.750 67.330 ;
        RECT 38.480 62.050 38.710 67.330 ;
        RECT 39.430 62.720 39.750 67.330 ;
        RECT 40.480 62.050 40.710 67.330 ;
        RECT 41.430 62.720 41.750 67.330 ;
        RECT 42.480 62.050 42.710 67.330 ;
        RECT 43.380 62.720 44.290 67.330 ;
        RECT 44.960 62.050 45.190 67.330 ;
        RECT 45.910 62.720 46.230 67.330 ;
        RECT 46.960 62.050 47.190 67.330 ;
        RECT 47.910 62.720 48.230 67.330 ;
        RECT 48.960 62.050 49.190 67.330 ;
        RECT 49.910 62.720 50.230 67.330 ;
        RECT 50.960 62.050 51.190 67.330 ;
        RECT 51.910 62.720 52.230 67.330 ;
        RECT 52.960 62.050 53.190 67.330 ;
        RECT 53.860 62.720 54.770 67.330 ;
        RECT 55.440 62.050 55.670 67.330 ;
        RECT 56.390 62.720 56.710 67.330 ;
        RECT 57.440 62.050 57.670 67.330 ;
        RECT 58.390 62.720 58.710 67.330 ;
        RECT 59.440 62.050 59.670 67.330 ;
        RECT 60.390 62.720 60.710 67.330 ;
        RECT 61.440 62.050 61.670 67.330 ;
        RECT 62.390 62.720 62.710 67.330 ;
        RECT 63.440 62.050 63.670 67.330 ;
        RECT 64.340 62.720 65.250 67.330 ;
        RECT 65.920 62.050 66.150 67.330 ;
        RECT 66.870 62.720 67.190 67.330 ;
        RECT 67.920 62.050 68.150 67.330 ;
        RECT 68.870 62.720 69.190 67.330 ;
        RECT 69.920 62.050 70.150 67.330 ;
        RECT 70.870 62.720 71.190 67.330 ;
        RECT 71.920 62.050 72.150 67.330 ;
        RECT 72.870 62.720 73.190 67.330 ;
        RECT 73.920 62.050 74.150 67.330 ;
        RECT 74.820 62.720 75.730 67.330 ;
        RECT 76.400 62.050 76.630 67.330 ;
        RECT 77.350 62.720 77.670 67.330 ;
        RECT 78.400 62.050 78.630 67.330 ;
        RECT 79.350 62.720 79.670 67.330 ;
        RECT 80.400 62.050 80.630 67.330 ;
        RECT 81.350 62.720 81.670 67.330 ;
        RECT 82.400 62.050 82.630 67.330 ;
        RECT 83.350 62.720 83.670 67.330 ;
        RECT 84.400 62.050 84.630 67.330 ;
        RECT 85.300 62.720 86.210 67.330 ;
        RECT 86.880 62.050 87.110 67.330 ;
        RECT 87.830 62.720 88.150 67.330 ;
        RECT 88.880 62.050 89.110 67.330 ;
        RECT 89.830 62.720 90.150 67.330 ;
        RECT 90.880 62.050 91.110 67.330 ;
        RECT 91.830 62.720 92.150 67.330 ;
        RECT 92.880 62.050 93.110 67.330 ;
        RECT 93.830 62.720 94.150 67.330 ;
        RECT 94.880 62.050 95.110 67.330 ;
        RECT 95.780 62.720 96.690 67.330 ;
        RECT 97.360 62.050 97.590 67.330 ;
        RECT 98.310 62.720 98.630 67.330 ;
        RECT 99.360 62.050 99.590 67.330 ;
        RECT 100.310 62.720 100.630 67.330 ;
        RECT 101.360 62.050 101.590 67.330 ;
        RECT 102.310 62.720 102.630 67.330 ;
        RECT 103.360 62.050 103.590 67.330 ;
        RECT 104.310 62.720 104.630 67.330 ;
        RECT 105.360 62.050 105.590 67.330 ;
        RECT 106.260 62.720 107.170 67.330 ;
        RECT 107.840 62.050 108.070 67.330 ;
        RECT 108.790 62.720 109.110 67.330 ;
        RECT 109.840 62.050 110.070 67.330 ;
        RECT 110.790 62.720 111.110 67.330 ;
        RECT 111.840 62.050 112.070 67.330 ;
        RECT 112.790 62.720 113.110 67.330 ;
        RECT 113.840 62.050 114.070 67.330 ;
        RECT 114.790 62.720 115.110 67.330 ;
        RECT 115.840 62.050 116.070 67.330 ;
        RECT 116.740 62.730 117.060 67.330 ;
        RECT 116.740 62.720 116.970 62.730 ;
        RECT 117.450 62.050 117.750 74.420 ;
        RECT 11.830 61.750 117.750 62.050 ;
        RECT 75.780 56.835 85.780 61.750 ;
        RECT 4.000 11.580 75.620 11.880 ;
        RECT 4.000 10.580 52.430 11.580 ;
        RECT 53.250 11.030 62.610 11.330 ;
        RECT 63.430 10.580 64.320 11.580 ;
        RECT 65.140 11.030 74.500 11.330 ;
        RECT 75.320 10.580 75.620 11.580 ;
        RECT 4.000 5.300 53.150 10.580 ;
        RECT 53.770 5.880 54.090 10.580 ;
        RECT 54.820 5.300 55.050 10.580 ;
        RECT 55.770 5.880 56.090 10.580 ;
        RECT 56.820 5.300 57.050 10.580 ;
        RECT 57.770 5.880 58.090 10.580 ;
        RECT 58.820 5.300 59.050 10.580 ;
        RECT 59.770 5.880 60.090 10.580 ;
        RECT 60.820 5.300 61.050 10.580 ;
        RECT 61.770 5.880 62.090 10.580 ;
        RECT 62.720 5.300 65.040 10.580 ;
        RECT 65.660 5.880 65.980 10.580 ;
        RECT 66.710 5.300 66.940 10.580 ;
        RECT 67.660 5.880 67.980 10.580 ;
        RECT 68.710 5.300 68.940 10.580 ;
        RECT 69.660 5.880 69.980 10.580 ;
        RECT 70.710 5.300 70.940 10.580 ;
        RECT 71.660 5.880 71.980 10.580 ;
        RECT 72.710 5.300 72.940 10.580 ;
        RECT 73.660 5.880 73.980 10.580 ;
        RECT 74.610 5.300 75.620 10.580 ;
        RECT 76.770 5.880 84.770 56.835 ;
        RECT 130.110 17.240 136.110 119.250 ;
        RECT 96.410 11.240 136.110 17.240 ;
        RECT 96.410 7.240 100.410 11.240 ;
        RECT 4.000 5.000 75.620 5.300 ;
      LAYER met2 ;
        RECT 4.000 5.000 6.000 220.760 ;
        RECT 7.000 5.000 9.000 220.760 ;
        RECT 120.850 171.200 140.580 171.900 ;
        RECT 30.990 113.800 40.990 133.020 ;
        RECT 119.660 130.100 120.460 170.800 ;
        RECT 120.850 130.100 121.850 171.200 ;
        RECT 107.050 120.800 121.850 130.100 ;
        RECT 125.450 120.800 126.450 171.200 ;
        RECT 130.050 120.800 131.050 171.200 ;
        RECT 134.650 120.800 135.650 171.200 ;
        RECT 139.580 120.800 140.580 171.200 ;
        RECT 140.970 121.190 141.770 170.800 ;
        RECT 107.050 120.100 140.580 120.800 ;
        RECT 107.050 113.800 117.050 120.100 ;
        RECT 12.560 112.800 117.050 113.800 ;
        RECT 12.560 112.030 12.880 112.800 ;
        RECT 14.460 112.030 14.780 112.800 ;
        RECT 16.460 112.030 16.780 112.800 ;
        RECT 18.460 112.030 18.780 112.800 ;
        RECT 20.460 112.030 20.780 112.800 ;
        RECT 22.410 112.030 23.320 112.800 ;
        RECT 24.940 112.030 25.260 112.800 ;
        RECT 26.940 112.030 27.260 112.800 ;
        RECT 28.940 112.030 29.260 112.800 ;
        RECT 30.940 112.030 31.260 112.800 ;
        RECT 32.890 112.030 33.800 112.800 ;
        RECT 35.420 112.030 35.740 112.800 ;
        RECT 37.420 112.030 37.740 112.800 ;
        RECT 39.420 112.030 39.740 112.800 ;
        RECT 41.420 112.030 41.740 112.800 ;
        RECT 43.370 112.030 44.280 112.800 ;
        RECT 45.900 112.030 46.220 112.800 ;
        RECT 47.900 112.030 48.220 112.800 ;
        RECT 49.900 112.030 50.220 112.800 ;
        RECT 51.900 112.030 52.220 112.800 ;
        RECT 53.850 112.030 54.760 112.800 ;
        RECT 56.380 112.030 56.700 112.800 ;
        RECT 58.380 112.030 58.700 112.800 ;
        RECT 60.380 112.030 60.700 112.800 ;
        RECT 62.380 112.030 62.700 112.800 ;
        RECT 64.330 112.030 65.240 112.800 ;
        RECT 66.860 112.030 67.180 112.800 ;
        RECT 68.860 112.030 69.180 112.800 ;
        RECT 70.860 112.030 71.180 112.800 ;
        RECT 72.860 112.030 73.180 112.800 ;
        RECT 74.810 112.030 75.720 112.800 ;
        RECT 77.340 112.030 77.660 112.800 ;
        RECT 79.340 112.030 79.660 112.800 ;
        RECT 81.340 112.030 81.660 112.800 ;
        RECT 83.340 112.030 83.660 112.800 ;
        RECT 85.290 112.030 86.200 112.800 ;
        RECT 87.820 112.030 88.140 112.800 ;
        RECT 89.820 112.030 90.140 112.800 ;
        RECT 91.820 112.030 92.140 112.800 ;
        RECT 93.820 112.030 94.140 112.800 ;
        RECT 95.770 112.030 96.680 112.800 ;
        RECT 98.300 112.030 98.620 112.800 ;
        RECT 100.300 112.030 100.620 112.800 ;
        RECT 102.300 112.030 102.620 112.800 ;
        RECT 104.300 112.030 104.620 112.800 ;
        RECT 106.250 112.030 107.160 112.800 ;
        RECT 108.780 112.030 109.100 112.800 ;
        RECT 110.780 112.030 111.100 112.800 ;
        RECT 112.780 112.030 113.100 112.800 ;
        RECT 114.780 112.030 115.100 112.800 ;
        RECT 116.730 112.030 117.050 112.800 ;
        RECT 12.560 111.030 117.050 112.030 ;
        RECT 12.560 110.190 12.880 111.030 ;
        RECT 14.460 110.190 14.780 111.030 ;
        RECT 16.460 110.190 16.780 111.030 ;
        RECT 18.460 110.190 18.780 111.030 ;
        RECT 20.460 110.190 20.780 111.030 ;
        RECT 22.410 110.190 23.320 111.030 ;
        RECT 24.940 110.190 25.260 111.030 ;
        RECT 26.940 110.190 27.260 111.030 ;
        RECT 28.940 110.190 29.260 111.030 ;
        RECT 30.940 110.190 31.260 111.030 ;
        RECT 32.890 110.190 33.800 111.030 ;
        RECT 35.420 110.190 35.740 111.030 ;
        RECT 37.420 110.190 37.740 111.030 ;
        RECT 39.420 110.190 39.740 111.030 ;
        RECT 41.420 110.190 41.740 111.030 ;
        RECT 43.370 110.190 44.280 111.030 ;
        RECT 45.900 110.190 46.220 111.030 ;
        RECT 47.900 110.190 48.220 111.030 ;
        RECT 49.900 110.190 50.220 111.030 ;
        RECT 51.900 110.190 52.220 111.030 ;
        RECT 53.850 110.190 54.760 111.030 ;
        RECT 56.380 110.190 56.700 111.030 ;
        RECT 58.380 110.190 58.700 111.030 ;
        RECT 60.380 110.190 60.700 111.030 ;
        RECT 62.380 110.190 62.700 111.030 ;
        RECT 64.330 110.190 65.240 111.030 ;
        RECT 66.860 110.190 67.180 111.030 ;
        RECT 68.860 110.190 69.180 111.030 ;
        RECT 70.860 110.190 71.180 111.030 ;
        RECT 72.860 110.190 73.180 111.030 ;
        RECT 74.810 110.190 75.720 111.030 ;
        RECT 77.340 110.190 77.660 111.030 ;
        RECT 79.340 110.190 79.660 111.030 ;
        RECT 81.340 110.190 81.660 111.030 ;
        RECT 83.340 110.190 83.660 111.030 ;
        RECT 85.290 110.190 86.200 111.030 ;
        RECT 87.820 110.190 88.140 111.030 ;
        RECT 89.820 110.190 90.140 111.030 ;
        RECT 91.820 110.190 92.140 111.030 ;
        RECT 93.820 110.190 94.140 111.030 ;
        RECT 95.770 110.190 96.680 111.030 ;
        RECT 98.300 110.190 98.620 111.030 ;
        RECT 100.300 110.190 100.620 111.030 ;
        RECT 102.300 110.190 102.620 111.030 ;
        RECT 104.300 110.190 104.620 111.030 ;
        RECT 106.250 110.190 107.160 111.030 ;
        RECT 108.780 110.190 109.100 111.030 ;
        RECT 110.780 110.190 111.100 111.030 ;
        RECT 112.780 110.190 113.100 111.030 ;
        RECT 114.780 110.190 115.100 111.030 ;
        RECT 116.730 110.190 117.050 111.030 ;
        RECT 12.530 109.190 117.050 110.190 ;
        RECT 12.530 107.380 14.530 109.190 ;
        RECT 14.950 107.830 20.350 108.740 ;
        RECT 20.650 107.380 22.650 109.190 ;
        RECT 23.010 107.380 25.010 109.190 ;
        RECT 25.430 107.830 30.830 108.740 ;
        RECT 31.130 107.380 33.130 109.190 ;
        RECT 33.490 107.380 35.490 109.190 ;
        RECT 35.910 107.830 41.310 108.740 ;
        RECT 41.610 107.380 43.610 109.190 ;
        RECT 43.970 107.380 45.970 109.190 ;
        RECT 46.390 107.830 51.790 108.740 ;
        RECT 52.090 107.380 54.090 109.190 ;
        RECT 54.450 107.380 56.450 109.190 ;
        RECT 56.870 107.830 62.270 108.740 ;
        RECT 62.570 107.380 64.570 109.190 ;
        RECT 64.930 107.380 66.930 109.190 ;
        RECT 67.350 107.830 72.750 108.740 ;
        RECT 73.050 107.380 75.050 109.190 ;
        RECT 75.410 107.380 77.410 109.190 ;
        RECT 77.830 107.830 83.230 108.740 ;
        RECT 83.530 107.380 85.530 109.190 ;
        RECT 85.890 107.380 87.890 109.190 ;
        RECT 88.310 107.830 93.710 108.740 ;
        RECT 94.010 107.380 96.010 109.190 ;
        RECT 96.370 107.380 98.370 109.190 ;
        RECT 98.790 107.830 104.190 108.740 ;
        RECT 104.490 107.380 106.490 109.190 ;
        RECT 106.850 107.380 108.850 109.190 ;
        RECT 109.270 107.830 114.670 108.740 ;
        RECT 114.970 107.380 116.970 109.190 ;
        RECT 12.530 106.380 117.060 107.380 ;
        RECT 12.570 105.540 12.890 106.380 ;
        RECT 14.470 105.540 14.790 106.380 ;
        RECT 16.470 105.540 16.790 106.380 ;
        RECT 18.470 105.540 18.790 106.380 ;
        RECT 20.470 105.540 20.790 106.380 ;
        RECT 22.420 105.540 23.330 106.380 ;
        RECT 24.950 105.540 25.270 106.380 ;
        RECT 26.950 105.540 27.270 106.380 ;
        RECT 28.950 105.540 29.270 106.380 ;
        RECT 30.950 105.540 31.270 106.380 ;
        RECT 32.900 105.540 33.810 106.380 ;
        RECT 35.430 105.540 35.750 106.380 ;
        RECT 37.430 105.540 37.750 106.380 ;
        RECT 39.430 105.540 39.750 106.380 ;
        RECT 41.430 105.540 41.750 106.380 ;
        RECT 43.380 105.540 44.290 106.380 ;
        RECT 45.910 105.540 46.230 106.380 ;
        RECT 47.910 105.540 48.230 106.380 ;
        RECT 49.910 105.540 50.230 106.380 ;
        RECT 51.910 105.540 52.230 106.380 ;
        RECT 53.860 105.540 54.770 106.380 ;
        RECT 56.390 105.540 56.710 106.380 ;
        RECT 58.390 105.540 58.710 106.380 ;
        RECT 60.390 105.540 60.710 106.380 ;
        RECT 62.390 105.540 62.710 106.380 ;
        RECT 64.340 105.540 65.250 106.380 ;
        RECT 66.870 105.540 67.190 106.380 ;
        RECT 68.870 105.540 69.190 106.380 ;
        RECT 70.870 105.540 71.190 106.380 ;
        RECT 72.870 105.540 73.190 106.380 ;
        RECT 74.820 105.540 75.730 106.380 ;
        RECT 77.350 105.540 77.670 106.380 ;
        RECT 79.350 105.540 79.670 106.380 ;
        RECT 81.350 105.540 81.670 106.380 ;
        RECT 83.350 105.540 83.670 106.380 ;
        RECT 85.300 105.540 86.210 106.380 ;
        RECT 87.830 105.540 88.150 106.380 ;
        RECT 89.830 105.540 90.150 106.380 ;
        RECT 91.830 105.540 92.150 106.380 ;
        RECT 93.830 105.540 94.150 106.380 ;
        RECT 95.780 105.540 96.690 106.380 ;
        RECT 98.310 105.540 98.630 106.380 ;
        RECT 100.310 105.540 100.630 106.380 ;
        RECT 102.310 105.540 102.630 106.380 ;
        RECT 104.310 105.540 104.630 106.380 ;
        RECT 106.260 105.540 107.170 106.380 ;
        RECT 108.790 105.540 109.110 106.380 ;
        RECT 110.790 105.540 111.110 106.380 ;
        RECT 112.790 105.540 113.110 106.380 ;
        RECT 114.790 105.540 115.110 106.380 ;
        RECT 116.740 105.540 117.060 106.380 ;
        RECT 12.530 104.540 117.060 105.540 ;
        RECT 12.570 103.770 12.890 104.540 ;
        RECT 14.470 103.770 14.790 104.540 ;
        RECT 16.470 103.770 16.790 104.540 ;
        RECT 18.470 103.770 18.790 104.540 ;
        RECT 20.470 103.770 20.790 104.540 ;
        RECT 22.420 103.770 23.330 104.540 ;
        RECT 24.950 103.770 25.270 104.540 ;
        RECT 26.950 103.770 27.270 104.540 ;
        RECT 28.950 103.770 29.270 104.540 ;
        RECT 30.950 103.770 31.270 104.540 ;
        RECT 32.900 103.770 33.810 104.540 ;
        RECT 35.430 103.770 35.750 104.540 ;
        RECT 37.430 103.770 37.750 104.540 ;
        RECT 39.430 103.770 39.750 104.540 ;
        RECT 41.430 103.770 41.750 104.540 ;
        RECT 43.380 103.770 44.290 104.540 ;
        RECT 45.910 103.770 46.230 104.540 ;
        RECT 47.910 103.770 48.230 104.540 ;
        RECT 49.910 103.770 50.230 104.540 ;
        RECT 51.910 103.770 52.230 104.540 ;
        RECT 53.860 103.770 54.770 104.540 ;
        RECT 56.390 103.770 56.710 104.540 ;
        RECT 58.390 103.770 58.710 104.540 ;
        RECT 60.390 103.770 60.710 104.540 ;
        RECT 62.390 103.770 62.710 104.540 ;
        RECT 64.340 103.770 65.250 104.540 ;
        RECT 66.870 103.770 67.190 104.540 ;
        RECT 68.870 103.770 69.190 104.540 ;
        RECT 70.870 103.770 71.190 104.540 ;
        RECT 72.870 103.770 73.190 104.540 ;
        RECT 74.820 103.770 75.730 104.540 ;
        RECT 77.350 103.770 77.670 104.540 ;
        RECT 79.350 103.770 79.670 104.540 ;
        RECT 81.350 103.770 81.670 104.540 ;
        RECT 83.350 103.770 83.670 104.540 ;
        RECT 85.300 103.770 86.210 104.540 ;
        RECT 87.830 103.770 88.150 104.540 ;
        RECT 89.830 103.770 90.150 104.540 ;
        RECT 91.830 103.770 92.150 104.540 ;
        RECT 93.830 103.770 94.150 104.540 ;
        RECT 95.780 103.770 96.690 104.540 ;
        RECT 98.310 103.770 98.630 104.540 ;
        RECT 100.310 103.770 100.630 104.540 ;
        RECT 102.310 103.770 102.630 104.540 ;
        RECT 104.310 103.770 104.630 104.540 ;
        RECT 106.260 103.770 107.170 104.540 ;
        RECT 108.790 103.770 109.110 104.540 ;
        RECT 110.790 103.770 111.110 104.540 ;
        RECT 112.790 103.770 113.110 104.540 ;
        RECT 114.790 103.770 115.110 104.540 ;
        RECT 116.740 103.770 117.060 104.540 ;
        RECT 12.530 100.450 117.060 103.770 ;
        RECT 12.560 99.450 117.050 100.450 ;
        RECT 12.560 98.680 12.880 99.450 ;
        RECT 14.460 98.680 14.780 99.450 ;
        RECT 16.460 98.680 16.780 99.450 ;
        RECT 18.460 98.680 18.780 99.450 ;
        RECT 20.460 98.680 20.780 99.450 ;
        RECT 22.410 98.680 23.320 99.450 ;
        RECT 24.940 98.680 25.260 99.450 ;
        RECT 26.940 98.680 27.260 99.450 ;
        RECT 28.940 98.680 29.260 99.450 ;
        RECT 30.940 98.680 31.260 99.450 ;
        RECT 32.890 98.680 33.800 99.450 ;
        RECT 35.420 98.680 35.740 99.450 ;
        RECT 37.420 98.680 37.740 99.450 ;
        RECT 39.420 98.680 39.740 99.450 ;
        RECT 41.420 98.680 41.740 99.450 ;
        RECT 43.370 98.680 44.280 99.450 ;
        RECT 45.900 98.680 46.220 99.450 ;
        RECT 47.900 98.680 48.220 99.450 ;
        RECT 49.900 98.680 50.220 99.450 ;
        RECT 51.900 98.680 52.220 99.450 ;
        RECT 53.850 98.680 54.760 99.450 ;
        RECT 56.380 98.680 56.700 99.450 ;
        RECT 58.380 98.680 58.700 99.450 ;
        RECT 60.380 98.680 60.700 99.450 ;
        RECT 62.380 98.680 62.700 99.450 ;
        RECT 64.330 98.680 65.240 99.450 ;
        RECT 66.860 98.680 67.180 99.450 ;
        RECT 68.860 98.680 69.180 99.450 ;
        RECT 70.860 98.680 71.180 99.450 ;
        RECT 72.860 98.680 73.180 99.450 ;
        RECT 74.810 98.680 75.720 99.450 ;
        RECT 77.340 98.680 77.660 99.450 ;
        RECT 79.340 98.680 79.660 99.450 ;
        RECT 81.340 98.680 81.660 99.450 ;
        RECT 83.340 98.680 83.660 99.450 ;
        RECT 85.290 98.680 86.200 99.450 ;
        RECT 87.820 98.680 88.140 99.450 ;
        RECT 89.820 98.680 90.140 99.450 ;
        RECT 91.820 98.680 92.140 99.450 ;
        RECT 93.820 98.680 94.140 99.450 ;
        RECT 95.770 98.680 96.680 99.450 ;
        RECT 98.300 98.680 98.620 99.450 ;
        RECT 100.300 98.680 100.620 99.450 ;
        RECT 102.300 98.680 102.620 99.450 ;
        RECT 104.300 98.680 104.620 99.450 ;
        RECT 106.250 98.680 107.160 99.450 ;
        RECT 108.780 98.680 109.100 99.450 ;
        RECT 110.780 98.680 111.100 99.450 ;
        RECT 112.780 98.680 113.100 99.450 ;
        RECT 114.780 98.680 115.100 99.450 ;
        RECT 116.730 98.680 117.050 99.450 ;
        RECT 12.560 97.680 117.050 98.680 ;
        RECT 12.560 96.840 12.880 97.680 ;
        RECT 14.460 96.840 14.780 97.680 ;
        RECT 16.460 96.840 16.780 97.680 ;
        RECT 18.460 96.840 18.780 97.680 ;
        RECT 20.460 96.840 20.780 97.680 ;
        RECT 22.410 96.840 23.320 97.680 ;
        RECT 24.940 96.840 25.260 97.680 ;
        RECT 26.940 96.840 27.260 97.680 ;
        RECT 28.940 96.840 29.260 97.680 ;
        RECT 30.940 96.840 31.260 97.680 ;
        RECT 32.890 96.840 33.800 97.680 ;
        RECT 35.420 96.840 35.740 97.680 ;
        RECT 37.420 96.840 37.740 97.680 ;
        RECT 39.420 96.840 39.740 97.680 ;
        RECT 41.420 96.840 41.740 97.680 ;
        RECT 43.370 96.840 44.280 97.680 ;
        RECT 45.900 96.840 46.220 97.680 ;
        RECT 47.900 96.840 48.220 97.680 ;
        RECT 49.900 96.840 50.220 97.680 ;
        RECT 51.900 96.840 52.220 97.680 ;
        RECT 53.850 96.840 54.760 97.680 ;
        RECT 56.380 96.840 56.700 97.680 ;
        RECT 58.380 96.840 58.700 97.680 ;
        RECT 60.380 96.840 60.700 97.680 ;
        RECT 62.380 96.840 62.700 97.680 ;
        RECT 64.330 96.840 65.240 97.680 ;
        RECT 66.860 96.840 67.180 97.680 ;
        RECT 68.860 96.840 69.180 97.680 ;
        RECT 70.860 96.840 71.180 97.680 ;
        RECT 72.860 96.840 73.180 97.680 ;
        RECT 74.810 96.840 75.720 97.680 ;
        RECT 77.340 96.840 77.660 97.680 ;
        RECT 79.340 96.840 79.660 97.680 ;
        RECT 81.340 96.840 81.660 97.680 ;
        RECT 83.340 96.840 83.660 97.680 ;
        RECT 85.290 96.840 86.200 97.680 ;
        RECT 87.820 96.840 88.140 97.680 ;
        RECT 89.820 96.840 90.140 97.680 ;
        RECT 91.820 96.840 92.140 97.680 ;
        RECT 93.820 96.840 94.140 97.680 ;
        RECT 95.770 96.840 96.680 97.680 ;
        RECT 98.300 96.840 98.620 97.680 ;
        RECT 100.300 96.840 100.620 97.680 ;
        RECT 102.300 96.840 102.620 97.680 ;
        RECT 104.300 96.840 104.620 97.680 ;
        RECT 106.250 96.840 107.160 97.680 ;
        RECT 108.780 96.840 109.100 97.680 ;
        RECT 110.780 96.840 111.100 97.680 ;
        RECT 112.780 96.840 113.100 97.680 ;
        RECT 114.780 96.840 115.100 97.680 ;
        RECT 116.730 96.840 117.050 97.680 ;
        RECT 12.530 95.840 117.050 96.840 ;
        RECT 12.530 94.030 14.530 95.840 ;
        RECT 14.950 94.480 20.350 95.390 ;
        RECT 20.650 94.030 22.650 95.840 ;
        RECT 23.010 94.030 25.010 95.840 ;
        RECT 25.430 94.480 30.830 95.390 ;
        RECT 31.130 94.030 33.130 95.840 ;
        RECT 33.490 94.030 35.490 95.840 ;
        RECT 35.910 94.480 41.310 95.390 ;
        RECT 41.610 94.030 43.610 95.840 ;
        RECT 43.970 94.030 45.970 95.840 ;
        RECT 46.390 94.480 51.790 95.390 ;
        RECT 52.090 94.030 54.090 95.840 ;
        RECT 54.450 94.030 56.450 95.840 ;
        RECT 56.870 94.480 62.270 95.390 ;
        RECT 62.570 94.030 64.570 95.840 ;
        RECT 64.930 94.030 66.930 95.840 ;
        RECT 67.350 94.480 72.750 95.390 ;
        RECT 73.050 94.030 75.050 95.840 ;
        RECT 75.410 94.030 77.410 95.840 ;
        RECT 77.830 94.480 83.230 95.390 ;
        RECT 83.530 94.030 85.530 95.840 ;
        RECT 85.890 94.030 87.890 95.840 ;
        RECT 88.310 94.480 93.710 95.390 ;
        RECT 94.010 94.030 96.010 95.840 ;
        RECT 96.370 94.030 98.370 95.840 ;
        RECT 98.790 94.480 104.190 95.390 ;
        RECT 104.490 94.030 106.490 95.840 ;
        RECT 106.850 94.030 108.850 95.840 ;
        RECT 109.270 94.480 114.670 95.390 ;
        RECT 114.970 94.030 116.970 95.840 ;
        RECT 12.530 93.030 117.060 94.030 ;
        RECT 12.570 92.190 12.890 93.030 ;
        RECT 14.470 92.190 14.790 93.030 ;
        RECT 16.470 92.190 16.790 93.030 ;
        RECT 18.470 92.190 18.790 93.030 ;
        RECT 20.470 92.190 20.790 93.030 ;
        RECT 22.420 92.190 23.330 93.030 ;
        RECT 24.950 92.190 25.270 93.030 ;
        RECT 26.950 92.190 27.270 93.030 ;
        RECT 28.950 92.190 29.270 93.030 ;
        RECT 30.950 92.190 31.270 93.030 ;
        RECT 32.900 92.190 33.810 93.030 ;
        RECT 35.430 92.190 35.750 93.030 ;
        RECT 37.430 92.190 37.750 93.030 ;
        RECT 39.430 92.190 39.750 93.030 ;
        RECT 41.430 92.190 41.750 93.030 ;
        RECT 43.380 92.190 44.290 93.030 ;
        RECT 45.910 92.190 46.230 93.030 ;
        RECT 47.910 92.190 48.230 93.030 ;
        RECT 49.910 92.190 50.230 93.030 ;
        RECT 51.910 92.190 52.230 93.030 ;
        RECT 53.860 92.190 54.770 93.030 ;
        RECT 56.390 92.190 56.710 93.030 ;
        RECT 58.390 92.190 58.710 93.030 ;
        RECT 60.390 92.190 60.710 93.030 ;
        RECT 62.390 92.190 62.710 93.030 ;
        RECT 64.340 92.190 65.250 93.030 ;
        RECT 66.870 92.190 67.190 93.030 ;
        RECT 68.870 92.190 69.190 93.030 ;
        RECT 70.870 92.190 71.190 93.030 ;
        RECT 72.870 92.190 73.190 93.030 ;
        RECT 74.820 92.190 75.730 93.030 ;
        RECT 77.350 92.190 77.670 93.030 ;
        RECT 79.350 92.190 79.670 93.030 ;
        RECT 81.350 92.190 81.670 93.030 ;
        RECT 83.350 92.190 83.670 93.030 ;
        RECT 85.300 92.190 86.210 93.030 ;
        RECT 87.830 92.190 88.150 93.030 ;
        RECT 89.830 92.190 90.150 93.030 ;
        RECT 91.830 92.190 92.150 93.030 ;
        RECT 93.830 92.190 94.150 93.030 ;
        RECT 95.780 92.190 96.690 93.030 ;
        RECT 98.310 92.190 98.630 93.030 ;
        RECT 100.310 92.190 100.630 93.030 ;
        RECT 102.310 92.190 102.630 93.030 ;
        RECT 104.310 92.190 104.630 93.030 ;
        RECT 106.260 92.190 107.170 93.030 ;
        RECT 108.790 92.190 109.110 93.030 ;
        RECT 110.790 92.190 111.110 93.030 ;
        RECT 112.790 92.190 113.110 93.030 ;
        RECT 114.790 92.190 115.110 93.030 ;
        RECT 116.740 92.190 117.060 93.030 ;
        RECT 12.530 91.420 117.060 92.190 ;
        RECT 9.520 91.190 117.060 91.420 ;
        RECT 9.520 90.420 12.890 91.190 ;
        RECT 14.470 90.420 14.790 91.190 ;
        RECT 16.470 90.420 16.790 91.190 ;
        RECT 18.470 90.420 18.790 91.190 ;
        RECT 20.470 90.420 20.790 91.190 ;
        RECT 22.420 90.420 23.330 91.190 ;
        RECT 24.950 90.420 25.270 91.190 ;
        RECT 26.950 90.420 27.270 91.190 ;
        RECT 28.950 90.420 29.270 91.190 ;
        RECT 30.950 90.420 31.270 91.190 ;
        RECT 32.900 90.420 33.810 91.190 ;
        RECT 35.430 90.420 35.750 91.190 ;
        RECT 37.430 90.420 37.750 91.190 ;
        RECT 39.430 90.420 39.750 91.190 ;
        RECT 41.430 90.420 41.750 91.190 ;
        RECT 43.380 90.420 44.290 91.190 ;
        RECT 45.910 90.420 46.230 91.190 ;
        RECT 47.910 90.420 48.230 91.190 ;
        RECT 49.910 90.420 50.230 91.190 ;
        RECT 51.910 90.420 52.230 91.190 ;
        RECT 53.860 90.420 54.770 91.190 ;
        RECT 56.390 90.420 56.710 91.190 ;
        RECT 58.390 90.420 58.710 91.190 ;
        RECT 60.390 90.420 60.710 91.190 ;
        RECT 62.390 90.420 62.710 91.190 ;
        RECT 64.340 90.420 65.250 91.190 ;
        RECT 66.870 90.420 67.190 91.190 ;
        RECT 68.870 90.420 69.190 91.190 ;
        RECT 70.870 90.420 71.190 91.190 ;
        RECT 72.870 90.420 73.190 91.190 ;
        RECT 74.820 90.420 75.730 91.190 ;
        RECT 77.350 90.420 77.670 91.190 ;
        RECT 79.350 90.420 79.670 91.190 ;
        RECT 81.350 90.420 81.670 91.190 ;
        RECT 83.350 90.420 83.670 91.190 ;
        RECT 85.300 90.420 86.210 91.190 ;
        RECT 87.830 90.420 88.150 91.190 ;
        RECT 89.830 90.420 90.150 91.190 ;
        RECT 91.830 90.420 92.150 91.190 ;
        RECT 93.830 90.420 94.150 91.190 ;
        RECT 95.780 90.420 96.690 91.190 ;
        RECT 98.310 90.420 98.630 91.190 ;
        RECT 100.310 90.420 100.630 91.190 ;
        RECT 102.310 90.420 102.630 91.190 ;
        RECT 104.310 90.420 104.630 91.190 ;
        RECT 106.260 90.420 107.170 91.190 ;
        RECT 108.790 90.420 109.110 91.190 ;
        RECT 110.790 90.420 111.110 91.190 ;
        RECT 112.790 90.420 113.110 91.190 ;
        RECT 114.790 90.420 115.110 91.190 ;
        RECT 116.740 90.420 117.060 91.190 ;
        RECT 9.520 89.430 117.060 90.420 ;
        RECT 9.520 89.420 116.970 89.430 ;
        RECT 9.520 82.580 11.520 89.420 ;
        RECT 118.380 87.100 120.380 93.930 ;
        RECT 12.560 86.100 120.380 87.100 ;
        RECT 12.560 85.330 12.880 86.100 ;
        RECT 14.460 85.330 14.780 86.100 ;
        RECT 16.460 85.330 16.780 86.100 ;
        RECT 18.460 85.330 18.780 86.100 ;
        RECT 20.460 85.330 20.780 86.100 ;
        RECT 22.410 85.330 23.320 86.100 ;
        RECT 24.940 85.330 25.260 86.100 ;
        RECT 26.940 85.330 27.260 86.100 ;
        RECT 28.940 85.330 29.260 86.100 ;
        RECT 30.940 85.330 31.260 86.100 ;
        RECT 32.890 85.330 33.800 86.100 ;
        RECT 35.420 85.330 35.740 86.100 ;
        RECT 37.420 85.330 37.740 86.100 ;
        RECT 39.420 85.330 39.740 86.100 ;
        RECT 41.420 85.330 41.740 86.100 ;
        RECT 43.370 85.330 44.280 86.100 ;
        RECT 45.900 85.330 46.220 86.100 ;
        RECT 47.900 85.330 48.220 86.100 ;
        RECT 49.900 85.330 50.220 86.100 ;
        RECT 51.900 85.330 52.220 86.100 ;
        RECT 53.850 85.330 54.760 86.100 ;
        RECT 56.380 85.330 56.700 86.100 ;
        RECT 58.380 85.330 58.700 86.100 ;
        RECT 60.380 85.330 60.700 86.100 ;
        RECT 62.380 85.330 62.700 86.100 ;
        RECT 64.330 85.330 65.240 86.100 ;
        RECT 66.860 85.330 67.180 86.100 ;
        RECT 68.860 85.330 69.180 86.100 ;
        RECT 70.860 85.330 71.180 86.100 ;
        RECT 72.860 85.330 73.180 86.100 ;
        RECT 74.810 85.330 75.720 86.100 ;
        RECT 77.340 85.330 77.660 86.100 ;
        RECT 79.340 85.330 79.660 86.100 ;
        RECT 81.340 85.330 81.660 86.100 ;
        RECT 83.340 85.330 83.660 86.100 ;
        RECT 85.290 85.330 86.200 86.100 ;
        RECT 87.820 85.330 88.140 86.100 ;
        RECT 89.820 85.330 90.140 86.100 ;
        RECT 91.820 85.330 92.140 86.100 ;
        RECT 93.820 85.330 94.140 86.100 ;
        RECT 95.770 85.330 96.680 86.100 ;
        RECT 98.300 85.330 98.620 86.100 ;
        RECT 100.300 85.330 100.620 86.100 ;
        RECT 102.300 85.330 102.620 86.100 ;
        RECT 104.300 85.330 104.620 86.100 ;
        RECT 106.250 85.330 107.160 86.100 ;
        RECT 108.780 85.330 109.100 86.100 ;
        RECT 110.780 85.330 111.100 86.100 ;
        RECT 112.780 85.330 113.100 86.100 ;
        RECT 114.780 85.330 115.100 86.100 ;
        RECT 116.730 85.330 120.380 86.100 ;
        RECT 12.560 85.100 120.380 85.330 ;
        RECT 12.560 84.330 117.050 85.100 ;
        RECT 12.560 83.490 12.880 84.330 ;
        RECT 14.460 83.490 14.780 84.330 ;
        RECT 16.460 83.490 16.780 84.330 ;
        RECT 18.460 83.490 18.780 84.330 ;
        RECT 20.460 83.490 20.780 84.330 ;
        RECT 22.410 83.490 23.320 84.330 ;
        RECT 24.940 83.490 25.260 84.330 ;
        RECT 26.940 83.490 27.260 84.330 ;
        RECT 28.940 83.490 29.260 84.330 ;
        RECT 30.940 83.490 31.260 84.330 ;
        RECT 32.890 83.490 33.800 84.330 ;
        RECT 35.420 83.490 35.740 84.330 ;
        RECT 37.420 83.490 37.740 84.330 ;
        RECT 39.420 83.490 39.740 84.330 ;
        RECT 41.420 83.490 41.740 84.330 ;
        RECT 43.370 83.490 44.280 84.330 ;
        RECT 45.900 83.490 46.220 84.330 ;
        RECT 47.900 83.490 48.220 84.330 ;
        RECT 49.900 83.490 50.220 84.330 ;
        RECT 51.900 83.490 52.220 84.330 ;
        RECT 53.850 83.490 54.760 84.330 ;
        RECT 56.380 83.490 56.700 84.330 ;
        RECT 58.380 83.490 58.700 84.330 ;
        RECT 60.380 83.490 60.700 84.330 ;
        RECT 62.380 83.490 62.700 84.330 ;
        RECT 64.330 83.490 65.240 84.330 ;
        RECT 66.860 83.490 67.180 84.330 ;
        RECT 68.860 83.490 69.180 84.330 ;
        RECT 70.860 83.490 71.180 84.330 ;
        RECT 72.860 83.490 73.180 84.330 ;
        RECT 74.810 83.490 75.720 84.330 ;
        RECT 77.340 83.490 77.660 84.330 ;
        RECT 79.340 83.490 79.660 84.330 ;
        RECT 81.340 83.490 81.660 84.330 ;
        RECT 83.340 83.490 83.660 84.330 ;
        RECT 85.290 83.490 86.200 84.330 ;
        RECT 87.820 83.490 88.140 84.330 ;
        RECT 89.820 83.490 90.140 84.330 ;
        RECT 91.820 83.490 92.140 84.330 ;
        RECT 93.820 83.490 94.140 84.330 ;
        RECT 95.770 83.490 96.680 84.330 ;
        RECT 98.300 83.490 98.620 84.330 ;
        RECT 100.300 83.490 100.620 84.330 ;
        RECT 102.300 83.490 102.620 84.330 ;
        RECT 104.300 83.490 104.620 84.330 ;
        RECT 106.250 83.490 107.160 84.330 ;
        RECT 108.780 83.490 109.100 84.330 ;
        RECT 110.780 83.490 111.100 84.330 ;
        RECT 112.780 83.490 113.100 84.330 ;
        RECT 114.780 83.490 115.100 84.330 ;
        RECT 116.730 83.490 117.050 84.330 ;
        RECT 12.530 82.490 117.050 83.490 ;
        RECT 12.530 80.680 14.530 82.490 ;
        RECT 14.950 81.130 20.350 82.040 ;
        RECT 20.650 80.680 22.650 82.490 ;
        RECT 23.010 80.680 25.010 82.490 ;
        RECT 25.430 81.130 30.830 82.040 ;
        RECT 31.130 80.680 33.130 82.490 ;
        RECT 33.490 80.680 35.490 82.490 ;
        RECT 35.910 81.130 41.310 82.040 ;
        RECT 41.610 80.680 43.610 82.490 ;
        RECT 43.970 80.680 45.970 82.490 ;
        RECT 46.390 81.130 51.790 82.040 ;
        RECT 52.090 80.680 54.090 82.490 ;
        RECT 54.450 80.680 56.450 82.490 ;
        RECT 56.870 81.130 62.270 82.040 ;
        RECT 62.570 80.680 64.570 82.490 ;
        RECT 64.930 80.680 66.930 82.490 ;
        RECT 67.350 81.130 72.750 82.040 ;
        RECT 73.050 80.680 75.050 82.490 ;
        RECT 75.410 80.680 77.410 82.490 ;
        RECT 77.830 81.130 83.230 82.040 ;
        RECT 83.530 80.680 85.530 82.490 ;
        RECT 85.890 80.680 87.890 82.490 ;
        RECT 88.310 81.130 93.710 82.040 ;
        RECT 94.010 80.680 96.010 82.490 ;
        RECT 96.370 80.680 98.370 82.490 ;
        RECT 98.790 81.130 104.190 82.040 ;
        RECT 104.490 80.680 106.490 82.490 ;
        RECT 106.850 80.680 108.850 82.490 ;
        RECT 109.270 81.130 114.670 82.040 ;
        RECT 114.970 80.680 116.970 82.490 ;
        RECT 12.530 79.680 117.060 80.680 ;
        RECT 12.570 78.840 12.890 79.680 ;
        RECT 14.470 78.840 14.790 79.680 ;
        RECT 16.470 78.840 16.790 79.680 ;
        RECT 18.470 78.840 18.790 79.680 ;
        RECT 20.470 78.840 20.790 79.680 ;
        RECT 22.420 78.840 23.330 79.680 ;
        RECT 24.950 78.840 25.270 79.680 ;
        RECT 26.950 78.840 27.270 79.680 ;
        RECT 28.950 78.840 29.270 79.680 ;
        RECT 30.950 78.840 31.270 79.680 ;
        RECT 32.900 78.840 33.810 79.680 ;
        RECT 35.430 78.840 35.750 79.680 ;
        RECT 37.430 78.840 37.750 79.680 ;
        RECT 39.430 78.840 39.750 79.680 ;
        RECT 41.430 78.840 41.750 79.680 ;
        RECT 43.380 78.840 44.290 79.680 ;
        RECT 45.910 78.840 46.230 79.680 ;
        RECT 47.910 78.840 48.230 79.680 ;
        RECT 49.910 78.840 50.230 79.680 ;
        RECT 51.910 78.840 52.230 79.680 ;
        RECT 53.860 78.840 54.770 79.680 ;
        RECT 56.390 78.840 56.710 79.680 ;
        RECT 58.390 78.840 58.710 79.680 ;
        RECT 60.390 78.840 60.710 79.680 ;
        RECT 62.390 78.840 62.710 79.680 ;
        RECT 64.340 78.840 65.250 79.680 ;
        RECT 66.870 78.840 67.190 79.680 ;
        RECT 68.870 78.840 69.190 79.680 ;
        RECT 70.870 78.840 71.190 79.680 ;
        RECT 72.870 78.840 73.190 79.680 ;
        RECT 74.820 78.840 75.730 79.680 ;
        RECT 77.350 78.840 77.670 79.680 ;
        RECT 79.350 78.840 79.670 79.680 ;
        RECT 81.350 78.840 81.670 79.680 ;
        RECT 83.350 78.840 83.670 79.680 ;
        RECT 85.300 78.840 86.210 79.680 ;
        RECT 87.830 78.840 88.150 79.680 ;
        RECT 89.830 78.840 90.150 79.680 ;
        RECT 91.830 78.840 92.150 79.680 ;
        RECT 93.830 78.840 94.150 79.680 ;
        RECT 95.780 78.840 96.690 79.680 ;
        RECT 98.310 78.840 98.630 79.680 ;
        RECT 100.310 78.840 100.630 79.680 ;
        RECT 102.310 78.840 102.630 79.680 ;
        RECT 104.310 78.840 104.630 79.680 ;
        RECT 106.260 78.840 107.170 79.680 ;
        RECT 108.790 78.840 109.110 79.680 ;
        RECT 110.790 78.840 111.110 79.680 ;
        RECT 112.790 78.840 113.110 79.680 ;
        RECT 114.790 78.840 115.110 79.680 ;
        RECT 116.740 78.840 117.060 79.680 ;
        RECT 12.530 77.840 117.060 78.840 ;
        RECT 12.570 77.070 12.890 77.840 ;
        RECT 14.470 77.070 14.790 77.840 ;
        RECT 16.470 77.070 16.790 77.840 ;
        RECT 18.470 77.070 18.790 77.840 ;
        RECT 20.470 77.070 20.790 77.840 ;
        RECT 22.420 77.070 23.330 77.840 ;
        RECT 24.950 77.070 25.270 77.840 ;
        RECT 26.950 77.070 27.270 77.840 ;
        RECT 28.950 77.070 29.270 77.840 ;
        RECT 30.950 77.070 31.270 77.840 ;
        RECT 32.900 77.070 33.810 77.840 ;
        RECT 35.430 77.070 35.750 77.840 ;
        RECT 37.430 77.070 37.750 77.840 ;
        RECT 39.430 77.070 39.750 77.840 ;
        RECT 41.430 77.070 41.750 77.840 ;
        RECT 43.380 77.070 44.290 77.840 ;
        RECT 45.910 77.070 46.230 77.840 ;
        RECT 47.910 77.070 48.230 77.840 ;
        RECT 49.910 77.070 50.230 77.840 ;
        RECT 51.910 77.070 52.230 77.840 ;
        RECT 53.860 77.070 54.770 77.840 ;
        RECT 56.390 77.070 56.710 77.840 ;
        RECT 58.390 77.070 58.710 77.840 ;
        RECT 60.390 77.070 60.710 77.840 ;
        RECT 62.390 77.070 62.710 77.840 ;
        RECT 64.340 77.070 65.250 77.840 ;
        RECT 66.870 77.070 67.190 77.840 ;
        RECT 68.870 77.070 69.190 77.840 ;
        RECT 70.870 77.070 71.190 77.840 ;
        RECT 72.870 77.070 73.190 77.840 ;
        RECT 74.820 77.070 75.730 77.840 ;
        RECT 77.350 77.070 77.670 77.840 ;
        RECT 79.350 77.070 79.670 77.840 ;
        RECT 81.350 77.070 81.670 77.840 ;
        RECT 83.350 77.070 83.670 77.840 ;
        RECT 85.300 77.070 86.210 77.840 ;
        RECT 87.830 77.070 88.150 77.840 ;
        RECT 89.830 77.070 90.150 77.840 ;
        RECT 91.830 77.070 92.150 77.840 ;
        RECT 93.830 77.070 94.150 77.840 ;
        RECT 95.780 77.070 96.690 77.840 ;
        RECT 98.310 77.070 98.630 77.840 ;
        RECT 100.310 77.070 100.630 77.840 ;
        RECT 102.310 77.070 102.630 77.840 ;
        RECT 104.310 77.070 104.630 77.840 ;
        RECT 106.260 77.070 107.170 77.840 ;
        RECT 108.790 77.070 109.110 77.840 ;
        RECT 110.790 77.070 111.110 77.840 ;
        RECT 112.790 77.070 113.110 77.840 ;
        RECT 114.790 77.070 115.110 77.840 ;
        RECT 116.740 77.070 117.060 77.840 ;
        RECT 12.530 73.750 117.060 77.070 ;
        RECT 12.560 72.750 117.050 73.750 ;
        RECT 12.560 71.980 12.880 72.750 ;
        RECT 14.460 71.980 14.780 72.750 ;
        RECT 16.460 71.980 16.780 72.750 ;
        RECT 18.460 71.980 18.780 72.750 ;
        RECT 20.460 71.980 20.780 72.750 ;
        RECT 22.410 71.980 23.320 72.750 ;
        RECT 24.940 71.980 25.260 72.750 ;
        RECT 26.940 71.980 27.260 72.750 ;
        RECT 28.940 71.980 29.260 72.750 ;
        RECT 30.940 71.980 31.260 72.750 ;
        RECT 32.890 71.980 33.800 72.750 ;
        RECT 35.420 71.980 35.740 72.750 ;
        RECT 37.420 71.980 37.740 72.750 ;
        RECT 39.420 71.980 39.740 72.750 ;
        RECT 41.420 71.980 41.740 72.750 ;
        RECT 43.370 71.980 44.280 72.750 ;
        RECT 45.900 71.980 46.220 72.750 ;
        RECT 47.900 71.980 48.220 72.750 ;
        RECT 49.900 71.980 50.220 72.750 ;
        RECT 51.900 71.980 52.220 72.750 ;
        RECT 53.850 71.980 54.760 72.750 ;
        RECT 56.380 71.980 56.700 72.750 ;
        RECT 58.380 71.980 58.700 72.750 ;
        RECT 60.380 71.980 60.700 72.750 ;
        RECT 62.380 71.980 62.700 72.750 ;
        RECT 64.330 71.980 65.240 72.750 ;
        RECT 66.860 71.980 67.180 72.750 ;
        RECT 68.860 71.980 69.180 72.750 ;
        RECT 70.860 71.980 71.180 72.750 ;
        RECT 72.860 71.980 73.180 72.750 ;
        RECT 74.810 71.980 75.720 72.750 ;
        RECT 77.340 71.980 77.660 72.750 ;
        RECT 79.340 71.980 79.660 72.750 ;
        RECT 81.340 71.980 81.660 72.750 ;
        RECT 83.340 71.980 83.660 72.750 ;
        RECT 85.290 71.980 86.200 72.750 ;
        RECT 87.820 71.980 88.140 72.750 ;
        RECT 89.820 71.980 90.140 72.750 ;
        RECT 91.820 71.980 92.140 72.750 ;
        RECT 93.820 71.980 94.140 72.750 ;
        RECT 95.770 71.980 96.680 72.750 ;
        RECT 98.300 71.980 98.620 72.750 ;
        RECT 100.300 71.980 100.620 72.750 ;
        RECT 102.300 71.980 102.620 72.750 ;
        RECT 104.300 71.980 104.620 72.750 ;
        RECT 106.250 71.980 107.160 72.750 ;
        RECT 108.780 71.980 109.100 72.750 ;
        RECT 110.780 71.980 111.100 72.750 ;
        RECT 112.780 71.980 113.100 72.750 ;
        RECT 114.780 71.980 115.100 72.750 ;
        RECT 116.730 71.980 117.050 72.750 ;
        RECT 12.560 70.980 117.050 71.980 ;
        RECT 12.560 70.140 12.880 70.980 ;
        RECT 14.460 70.140 14.780 70.980 ;
        RECT 16.460 70.140 16.780 70.980 ;
        RECT 18.460 70.140 18.780 70.980 ;
        RECT 20.460 70.140 20.780 70.980 ;
        RECT 22.410 70.140 23.320 70.980 ;
        RECT 24.940 70.140 25.260 70.980 ;
        RECT 26.940 70.140 27.260 70.980 ;
        RECT 28.940 70.140 29.260 70.980 ;
        RECT 30.940 70.140 31.260 70.980 ;
        RECT 32.890 70.140 33.800 70.980 ;
        RECT 35.420 70.140 35.740 70.980 ;
        RECT 37.420 70.140 37.740 70.980 ;
        RECT 39.420 70.140 39.740 70.980 ;
        RECT 41.420 70.140 41.740 70.980 ;
        RECT 43.370 70.140 44.280 70.980 ;
        RECT 45.900 70.140 46.220 70.980 ;
        RECT 47.900 70.140 48.220 70.980 ;
        RECT 49.900 70.140 50.220 70.980 ;
        RECT 51.900 70.140 52.220 70.980 ;
        RECT 53.850 70.140 54.760 70.980 ;
        RECT 56.380 70.140 56.700 70.980 ;
        RECT 58.380 70.140 58.700 70.980 ;
        RECT 60.380 70.140 60.700 70.980 ;
        RECT 62.380 70.140 62.700 70.980 ;
        RECT 64.330 70.140 65.240 70.980 ;
        RECT 66.860 70.140 67.180 70.980 ;
        RECT 68.860 70.140 69.180 70.980 ;
        RECT 70.860 70.140 71.180 70.980 ;
        RECT 72.860 70.140 73.180 70.980 ;
        RECT 74.810 70.140 75.720 70.980 ;
        RECT 77.340 70.140 77.660 70.980 ;
        RECT 79.340 70.140 79.660 70.980 ;
        RECT 81.340 70.140 81.660 70.980 ;
        RECT 83.340 70.140 83.660 70.980 ;
        RECT 85.290 70.140 86.200 70.980 ;
        RECT 87.820 70.140 88.140 70.980 ;
        RECT 89.820 70.140 90.140 70.980 ;
        RECT 91.820 70.140 92.140 70.980 ;
        RECT 93.820 70.140 94.140 70.980 ;
        RECT 95.770 70.140 96.680 70.980 ;
        RECT 98.300 70.140 98.620 70.980 ;
        RECT 100.300 70.140 100.620 70.980 ;
        RECT 102.300 70.140 102.620 70.980 ;
        RECT 104.300 70.140 104.620 70.980 ;
        RECT 106.250 70.140 107.160 70.980 ;
        RECT 108.780 70.140 109.100 70.980 ;
        RECT 110.780 70.140 111.100 70.980 ;
        RECT 112.780 70.140 113.100 70.980 ;
        RECT 114.780 70.140 115.100 70.980 ;
        RECT 116.730 70.140 117.050 70.980 ;
        RECT 12.530 69.140 117.050 70.140 ;
        RECT 12.530 67.330 14.530 69.140 ;
        RECT 14.950 67.780 20.350 68.690 ;
        RECT 20.650 67.330 22.650 69.140 ;
        RECT 23.010 67.330 25.010 69.140 ;
        RECT 25.430 67.780 30.830 68.690 ;
        RECT 31.130 67.330 33.130 69.140 ;
        RECT 33.490 67.330 35.490 69.140 ;
        RECT 35.910 67.780 41.310 68.690 ;
        RECT 41.610 67.330 43.610 69.140 ;
        RECT 43.970 67.330 45.970 69.140 ;
        RECT 46.390 67.780 51.790 68.690 ;
        RECT 52.090 67.330 54.090 69.140 ;
        RECT 54.450 67.330 56.450 69.140 ;
        RECT 56.870 67.780 62.270 68.690 ;
        RECT 62.570 67.330 64.570 69.140 ;
        RECT 64.930 67.330 66.930 69.140 ;
        RECT 67.350 67.780 72.750 68.690 ;
        RECT 73.050 67.330 75.050 69.140 ;
        RECT 75.410 67.330 77.410 69.140 ;
        RECT 77.830 67.780 83.230 68.690 ;
        RECT 83.530 67.330 85.530 69.140 ;
        RECT 85.890 67.330 87.890 69.140 ;
        RECT 88.310 67.780 93.710 68.690 ;
        RECT 94.010 67.330 96.010 69.140 ;
        RECT 96.370 67.330 98.370 69.140 ;
        RECT 98.790 67.780 104.190 68.690 ;
        RECT 104.490 67.330 106.490 69.140 ;
        RECT 106.850 67.330 108.850 69.140 ;
        RECT 109.270 67.780 114.670 68.690 ;
        RECT 114.970 67.330 116.970 69.140 ;
        RECT 12.530 66.330 117.060 67.330 ;
        RECT 12.570 65.490 12.890 66.330 ;
        RECT 14.470 65.490 14.790 66.330 ;
        RECT 16.470 65.490 16.790 66.330 ;
        RECT 18.470 65.490 18.790 66.330 ;
        RECT 20.470 65.490 20.790 66.330 ;
        RECT 22.420 65.490 23.330 66.330 ;
        RECT 24.950 65.490 25.270 66.330 ;
        RECT 26.950 65.490 27.270 66.330 ;
        RECT 28.950 65.490 29.270 66.330 ;
        RECT 30.950 65.490 31.270 66.330 ;
        RECT 32.900 65.490 33.810 66.330 ;
        RECT 35.430 65.490 35.750 66.330 ;
        RECT 37.430 65.490 37.750 66.330 ;
        RECT 39.430 65.490 39.750 66.330 ;
        RECT 41.430 65.490 41.750 66.330 ;
        RECT 43.380 65.490 44.290 66.330 ;
        RECT 45.910 65.490 46.230 66.330 ;
        RECT 47.910 65.490 48.230 66.330 ;
        RECT 49.910 65.490 50.230 66.330 ;
        RECT 51.910 65.490 52.230 66.330 ;
        RECT 53.860 65.490 54.770 66.330 ;
        RECT 56.390 65.490 56.710 66.330 ;
        RECT 58.390 65.490 58.710 66.330 ;
        RECT 60.390 65.490 60.710 66.330 ;
        RECT 62.390 65.490 62.710 66.330 ;
        RECT 64.340 65.490 65.250 66.330 ;
        RECT 66.870 65.490 67.190 66.330 ;
        RECT 68.870 65.490 69.190 66.330 ;
        RECT 70.870 65.490 71.190 66.330 ;
        RECT 72.870 65.490 73.190 66.330 ;
        RECT 74.820 65.490 75.730 66.330 ;
        RECT 77.350 65.490 77.670 66.330 ;
        RECT 79.350 65.490 79.670 66.330 ;
        RECT 81.350 65.490 81.670 66.330 ;
        RECT 83.350 65.490 83.670 66.330 ;
        RECT 85.300 65.490 86.210 66.330 ;
        RECT 87.830 65.490 88.150 66.330 ;
        RECT 89.830 65.490 90.150 66.330 ;
        RECT 91.830 65.490 92.150 66.330 ;
        RECT 93.830 65.490 94.150 66.330 ;
        RECT 95.780 65.490 96.690 66.330 ;
        RECT 98.310 65.490 98.630 66.330 ;
        RECT 100.310 65.490 100.630 66.330 ;
        RECT 102.310 65.490 102.630 66.330 ;
        RECT 104.310 65.490 104.630 66.330 ;
        RECT 106.260 65.490 107.170 66.330 ;
        RECT 108.790 65.490 109.110 66.330 ;
        RECT 110.790 65.490 111.110 66.330 ;
        RECT 112.790 65.490 113.110 66.330 ;
        RECT 114.790 65.490 115.110 66.330 ;
        RECT 116.740 65.490 117.060 66.330 ;
        RECT 12.530 64.490 117.060 65.490 ;
        RECT 12.570 63.720 12.890 64.490 ;
        RECT 14.470 63.720 14.790 64.490 ;
        RECT 16.470 63.720 16.790 64.490 ;
        RECT 18.470 63.720 18.790 64.490 ;
        RECT 20.470 63.720 20.790 64.490 ;
        RECT 22.420 63.720 23.330 64.490 ;
        RECT 24.950 63.720 25.270 64.490 ;
        RECT 26.950 63.720 27.270 64.490 ;
        RECT 28.950 63.720 29.270 64.490 ;
        RECT 30.950 63.720 31.270 64.490 ;
        RECT 32.900 63.720 33.810 64.490 ;
        RECT 35.430 63.720 35.750 64.490 ;
        RECT 37.430 63.720 37.750 64.490 ;
        RECT 39.430 63.720 39.750 64.490 ;
        RECT 41.430 63.720 41.750 64.490 ;
        RECT 43.380 63.720 44.290 64.490 ;
        RECT 45.910 63.720 46.230 64.490 ;
        RECT 47.910 63.720 48.230 64.490 ;
        RECT 49.910 63.720 50.230 64.490 ;
        RECT 51.910 63.720 52.230 64.490 ;
        RECT 53.860 63.720 54.770 64.490 ;
        RECT 56.390 63.720 56.710 64.490 ;
        RECT 58.390 63.720 58.710 64.490 ;
        RECT 60.390 63.720 60.710 64.490 ;
        RECT 62.390 63.720 62.710 64.490 ;
        RECT 64.340 63.720 65.250 64.490 ;
        RECT 66.870 63.720 67.190 64.490 ;
        RECT 68.870 63.720 69.190 64.490 ;
        RECT 70.870 63.720 71.190 64.490 ;
        RECT 72.870 63.720 73.190 64.490 ;
        RECT 74.820 63.720 75.730 64.490 ;
        RECT 77.350 63.720 77.670 64.490 ;
        RECT 79.350 63.720 79.670 64.490 ;
        RECT 81.350 63.720 81.670 64.490 ;
        RECT 83.350 63.720 83.670 64.490 ;
        RECT 85.300 63.720 86.210 64.490 ;
        RECT 87.830 63.720 88.150 64.490 ;
        RECT 89.830 63.720 90.150 64.490 ;
        RECT 91.830 63.720 92.150 64.490 ;
        RECT 93.830 63.720 94.150 64.490 ;
        RECT 95.780 63.720 96.690 64.490 ;
        RECT 98.310 63.720 98.630 64.490 ;
        RECT 100.310 63.720 100.630 64.490 ;
        RECT 102.310 63.720 102.630 64.490 ;
        RECT 104.310 63.720 104.630 64.490 ;
        RECT 106.260 63.720 107.170 64.490 ;
        RECT 108.790 63.720 109.110 64.490 ;
        RECT 110.790 63.720 111.110 64.490 ;
        RECT 112.790 63.720 113.110 64.490 ;
        RECT 114.790 63.720 115.110 64.490 ;
        RECT 116.740 63.720 117.060 64.490 ;
        RECT 12.530 62.730 117.060 63.720 ;
        RECT 12.530 62.720 116.970 62.730 ;
        RECT 136.580 17.240 140.580 120.100 ;
        RECT 53.250 11.030 74.500 11.330 ;
        RECT 53.770 9.580 62.090 11.030 ;
        RECT 53.770 8.740 54.090 9.580 ;
        RECT 55.770 8.740 56.090 9.580 ;
        RECT 57.770 8.740 58.090 9.580 ;
        RECT 59.770 8.740 60.090 9.580 ;
        RECT 61.770 8.740 62.090 9.580 ;
        RECT 53.770 7.740 62.090 8.740 ;
        RECT 53.770 6.880 54.090 7.740 ;
        RECT 55.770 6.880 56.090 7.740 ;
        RECT 57.770 6.880 58.090 7.740 ;
        RECT 59.770 6.880 60.090 7.740 ;
        RECT 61.770 6.880 62.090 7.740 ;
        RECT 53.770 5.880 62.090 6.880 ;
        RECT 65.660 9.580 84.770 10.580 ;
        RECT 65.660 8.710 65.980 9.580 ;
        RECT 67.660 8.710 67.980 9.580 ;
        RECT 69.660 8.710 69.980 9.580 ;
        RECT 71.660 8.710 71.980 9.580 ;
        RECT 73.660 8.710 84.770 9.580 ;
        RECT 65.660 7.710 84.770 8.710 ;
        RECT 65.660 6.880 65.980 7.710 ;
        RECT 67.660 6.880 67.980 7.710 ;
        RECT 69.660 6.880 69.980 7.710 ;
        RECT 71.660 6.880 71.980 7.710 ;
        RECT 73.660 6.880 84.770 7.710 ;
        RECT 96.410 7.240 100.410 17.240 ;
        RECT 134.910 13.240 140.580 17.240 ;
        RECT 134.910 7.240 138.910 13.240 ;
        RECT 65.660 5.880 84.770 6.880 ;
        RECT 60.090 4.170 62.090 5.880 ;
        RECT 60.090 2.170 79.720 4.170 ;
        RECT 77.720 1.570 79.720 2.170 ;
      LAYER met3 ;
        RECT 125.130 223.860 126.030 224.760 ;
        RECT 127.870 223.860 128.770 224.760 ;
        RECT 130.630 223.860 131.530 224.760 ;
        RECT 1.000 5.000 3.000 220.760 ;
        RECT 4.000 5.000 6.000 220.760 ;
        RECT 7.000 173.370 9.000 220.760 ;
        RECT 14.000 219.000 114.000 221.000 ;
        RECT 59.000 196.000 64.000 198.000 ;
        RECT 62.000 194.000 64.000 196.000 ;
        RECT 62.000 192.000 67.000 194.000 ;
        RECT 59.000 188.000 64.000 190.000 ;
        RECT 62.000 186.000 64.000 188.000 ;
        RECT 62.000 184.000 67.000 186.000 ;
        RECT 61.980 173.370 63.980 178.370 ;
        RECT 7.000 168.370 63.980 173.370 ;
        RECT 119.660 169.800 141.770 170.800 ;
        RECT 7.000 5.000 9.000 168.370 ;
        RECT 119.660 163.800 120.460 169.800 ;
        RECT 140.970 163.800 141.770 169.800 ;
        RECT 119.660 162.800 141.770 163.800 ;
        RECT 62.000 158.000 67.000 160.000 ;
        RECT 62.000 156.000 64.000 158.000 ;
        RECT 59.000 154.000 64.000 156.000 ;
        RECT 119.660 156.800 120.460 162.800 ;
        RECT 140.970 156.800 141.770 162.800 ;
        RECT 119.660 155.800 141.770 156.800 ;
        RECT 62.000 150.000 67.000 152.000 ;
        RECT 62.000 148.000 64.000 150.000 ;
        RECT 59.000 146.000 64.000 148.000 ;
        RECT 119.660 149.800 120.460 155.800 ;
        RECT 140.970 149.800 141.770 155.800 ;
        RECT 119.660 148.800 141.770 149.800 ;
        RECT 119.660 142.800 120.460 148.800 ;
        RECT 140.970 142.800 141.770 148.800 ;
        RECT 119.660 141.800 141.770 142.800 ;
        RECT 119.660 135.800 120.460 141.800 ;
        RECT 140.970 135.800 141.770 141.800 ;
        RECT 119.660 134.800 141.770 135.800 ;
        RECT 30.990 123.020 40.990 133.020 ;
        RECT 119.660 133.000 120.460 134.800 ;
        RECT 89.000 128.800 120.460 133.000 ;
        RECT 140.970 128.800 141.770 134.800 ;
        RECT 89.000 127.800 141.770 128.800 ;
        RECT 89.000 124.780 120.460 127.800 ;
        RECT 140.970 124.780 141.770 127.800 ;
        RECT 89.000 123.000 141.770 124.780 ;
        RECT 119.660 121.190 141.770 123.000 ;
        RECT 9.520 108.740 12.160 109.290 ;
        RECT 119.660 109.280 129.660 121.190 ;
        RECT 117.830 108.740 129.660 109.280 ;
        RECT 9.520 107.830 129.660 108.740 ;
        RECT 9.520 107.290 12.160 107.830 ;
        RECT 9.520 95.940 11.520 107.290 ;
        RECT 117.830 107.280 129.660 107.830 ;
        RECT 118.380 100.360 129.660 107.280 ;
        RECT 9.520 95.390 12.070 95.940 ;
        RECT 118.380 95.930 120.380 100.360 ;
        RECT 117.740 95.390 120.380 95.930 ;
        RECT 9.520 94.480 120.380 95.390 ;
        RECT 9.520 93.940 12.070 94.480 ;
        RECT 117.740 93.930 120.380 94.480 ;
        RECT 9.520 82.580 11.520 88.580 ;
        RECT 118.380 87.930 120.380 93.930 ;
        RECT 9.520 82.040 12.160 82.580 ;
        RECT 117.830 82.040 120.380 82.580 ;
        RECT 9.520 81.130 120.380 82.040 ;
        RECT 9.520 80.580 12.160 81.130 ;
        RECT 117.830 80.580 120.380 81.130 ;
        RECT 9.520 69.230 11.520 80.580 ;
        RECT 118.380 69.230 120.380 80.580 ;
        RECT 9.520 68.690 12.070 69.230 ;
        RECT 117.740 68.690 120.380 69.230 ;
        RECT 9.520 67.780 120.380 68.690 ;
        RECT 9.520 67.230 12.070 67.780 ;
        RECT 117.740 67.230 120.380 67.780 ;
        RECT 125.660 21.240 129.660 100.360 ;
        RECT 115.510 17.240 129.660 21.240 ;
        RECT 96.410 7.240 100.410 17.240 ;
        RECT 115.510 7.230 119.510 17.240 ;
        RECT 134.910 7.240 138.910 17.240 ;
        RECT 0.930 1.000 1.830 1.900 ;
        RECT 20.250 1.000 21.150 1.900 ;
        RECT 39.570 1.000 40.470 1.900 ;
        RECT 58.890 1.000 59.790 1.900 ;
        RECT 77.720 1.570 79.720 4.170 ;
      LAYER met4 ;
        RECT 15.030 223.960 15.330 224.760 ;
        RECT 17.790 223.960 18.090 224.760 ;
        RECT 20.550 223.960 20.850 224.760 ;
        RECT 23.310 223.960 23.610 224.760 ;
        RECT 26.070 223.960 26.370 224.760 ;
        RECT 28.830 223.960 29.130 224.760 ;
        RECT 31.590 223.960 31.890 224.760 ;
        RECT 34.350 223.960 34.650 224.760 ;
        RECT 37.110 223.960 37.410 224.760 ;
        RECT 39.870 223.960 40.170 224.760 ;
        RECT 42.630 223.960 42.930 224.760 ;
        RECT 45.390 223.960 45.690 224.760 ;
        RECT 48.150 223.960 48.450 224.760 ;
        RECT 50.910 223.960 51.210 224.760 ;
        RECT 53.670 223.960 53.970 224.760 ;
        RECT 56.430 223.960 56.730 224.760 ;
        RECT 59.190 223.960 59.490 224.760 ;
        RECT 61.950 223.960 62.250 224.760 ;
        RECT 64.710 223.960 65.010 224.760 ;
        RECT 67.470 223.960 67.770 224.760 ;
        RECT 70.230 223.960 70.530 224.760 ;
        RECT 72.990 223.960 73.290 224.760 ;
        RECT 75.750 223.960 76.050 224.760 ;
        RECT 78.510 223.960 78.810 224.760 ;
        RECT 81.270 223.960 81.570 224.760 ;
        RECT 84.030 223.960 84.330 224.760 ;
        RECT 86.790 223.960 87.090 224.760 ;
        RECT 89.550 223.960 89.850 224.760 ;
        RECT 92.310 223.960 92.610 224.760 ;
        RECT 95.070 223.960 95.370 224.760 ;
        RECT 97.830 223.960 98.130 224.760 ;
        RECT 100.590 223.960 100.890 224.760 ;
        RECT 103.350 223.960 103.650 224.760 ;
        RECT 106.110 223.960 106.410 224.760 ;
        RECT 108.870 223.960 109.170 224.760 ;
        RECT 111.630 223.960 111.930 224.760 ;
        RECT 114.390 223.960 114.690 224.760 ;
        RECT 117.150 223.960 117.450 224.760 ;
        RECT 119.910 223.960 120.210 224.760 ;
        RECT 122.670 223.960 122.970 224.760 ;
        RECT 4.800 223.660 122.970 223.960 ;
        RECT 125.130 223.860 126.030 224.760 ;
        RECT 127.870 223.860 128.770 224.760 ;
        RECT 130.630 223.860 131.530 224.760 ;
        RECT 4.800 220.760 5.100 223.660 ;
        RECT 34.350 223.610 34.650 223.660 ;
        RECT 39.870 223.580 40.170 223.660 ;
        RECT 12.000 219.000 114.000 221.000 ;
        RECT 12.000 121.000 14.000 219.000 ;
        RECT 35.000 196.000 61.000 198.000 ;
        RECT 62.000 196.000 91.000 198.000 ;
        RECT 35.000 133.020 37.000 196.000 ;
        RECT 62.000 194.000 64.000 196.000 ;
        RECT 39.000 192.000 64.000 194.000 ;
        RECT 65.000 192.000 87.000 194.000 ;
        RECT 39.000 148.000 41.000 192.000 ;
        RECT 43.000 188.000 61.000 190.000 ;
        RECT 62.000 188.000 83.000 190.000 ;
        RECT 43.000 152.000 45.000 188.000 ;
        RECT 62.000 186.000 64.000 188.000 ;
        RECT 47.000 184.000 64.000 186.000 ;
        RECT 65.000 184.000 79.000 186.000 ;
        RECT 47.000 156.000 49.000 184.000 ;
        RECT 51.000 180.000 75.000 182.000 ;
        RECT 51.000 160.000 53.000 180.000 ;
        RECT 62.000 178.370 64.000 180.000 ;
        RECT 61.980 171.000 64.000 178.370 ;
        RECT 61.980 168.370 63.980 171.000 ;
        RECT 73.000 160.000 75.000 180.000 ;
        RECT 51.000 158.000 64.000 160.000 ;
        RECT 65.000 158.000 75.000 160.000 ;
        RECT 62.000 156.000 64.000 158.000 ;
        RECT 77.000 156.000 79.000 184.000 ;
        RECT 47.000 154.000 61.000 156.000 ;
        RECT 62.000 154.000 79.000 156.000 ;
        RECT 81.000 152.000 83.000 188.000 ;
        RECT 43.000 150.000 64.000 152.000 ;
        RECT 65.000 150.000 83.000 152.000 ;
        RECT 62.000 148.000 64.000 150.000 ;
        RECT 85.000 148.000 87.000 192.000 ;
        RECT 39.000 146.000 61.000 148.000 ;
        RECT 62.000 146.000 87.000 148.000 ;
        RECT 30.990 123.020 40.990 133.020 ;
        RECT 89.000 123.000 91.000 196.000 ;
        RECT 112.000 121.000 114.000 219.000 ;
        RECT 12.000 119.000 114.000 121.000 ;
        RECT 96.410 7.240 100.410 17.240 ;
        RECT 0.930 1.000 1.830 1.900 ;
        RECT 20.250 1.000 21.150 1.900 ;
        RECT 39.570 1.000 40.470 1.900 ;
        RECT 58.890 1.000 59.790 1.900 ;
        RECT 77.720 1.570 79.720 4.170 ;
        RECT 97.230 1.575 98.705 7.240 ;
        RECT 115.510 7.230 119.510 17.230 ;
        RECT 134.910 7.240 138.910 17.240 ;
        RECT 116.550 1.575 118.025 7.230 ;
        RECT 135.870 1.575 137.345 7.240 ;
        RECT 78.210 1.000 79.110 1.570 ;
        RECT 97.530 1.000 98.430 1.575 ;
        RECT 116.850 1.000 117.750 1.575 ;
        RECT 136.170 1.000 137.070 1.575 ;
  END
END tt_um_noritsuna_Vctrl_LC_oscillator
END LIBRARY

